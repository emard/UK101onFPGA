library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity rom_bas is
	port (
		clk: in std_logic;
		addr: in std_logic_vector(12 downto 0);
		data: out std_logic_vector(7 downto 0)
	);
end entity;

architecture Behavioral of rom_bas is
	type romDef is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant romData: romDef := (
x"39", x"C6", x"55", x"C5", x"3F", x"CA", x"0B", x"C7",
x"22", x"C9", x"00", x"CD", x"4E", x"C9", x"98", x"DE",
x"B8", x"C6", x"90", x"C6", x"3B", x"C7", x"19", x"C6",
x"9B", x"C6", x"E5", x"C6", x"4E", x"C7", x"37", x"C6",
x"5E", x"C7", x"80", x"DE", x"8C", x"DE", x"26", x"F2",
x"F4", x"F0", x"DD", x"CF", x"28", x"D4", x"2E", x"C8",
x"60", x"C6", x"B4", x"C4", x"8B", x"C6", x"60", x"C4",
x"D8", x"D7", x"62", x"D8", x"F5", x"D7", x"0A", x"00",
x"AD", x"CF", x"CE", x"CF", x"AC", x"DA", x"C0", x"DB",
x"BD", x"D5", x"1B", x"DB", x"FC", x"DB", x"03", x"DC",
x"4C", x"DC", x"99", x"DC", x"1E", x"D4", x"8C", x"D3",
x"8C", x"D0", x"BD", x"D3", x"9B", x"D3", x"FC", x"D2",
x"10", x"D3", x"3C", x"D3", x"47", x"D3", x"79", x"6E",
x"D4", x"79", x"57", x"D4", x"7B", x"FD", x"D5", x"7B",
x"CC", x"D6", x"7F", x"B5", x"DA", x"50", x"68", x"CC",
x"46", x"65", x"CC", x"7D", x"EE", x"DA", x"5A", x"D7",
x"CB", x"64", x"95", x"CC", x"45", x"4E", x"C4", x"46",
x"4F", x"D2", x"4E", x"45", x"58", x"D4", x"44", x"41",
x"54", x"C1", x"49", x"4E", x"50", x"55", x"D4", x"44",
x"49", x"CD", x"52", x"45", x"41", x"C4", x"4D", x"4F",
x"D6", x"47", x"4F", x"54", x"CF", x"52", x"55", x"CE",
x"49", x"C6", x"52", x"45", x"53", x"54", x"4F", x"52",
x"C5", x"47", x"4F", x"53", x"55", x"C2", x"52", x"45",
x"54", x"55", x"52", x"CE", x"52", x"45", x"CD", x"53",
x"54", x"4F", x"D0", x"4F", x"CE", x"44", x"52", x"41",
x"D7", x"50", x"4C", x"4F", x"D4", x"4C", x"4F", x"41",
x"C4", x"53", x"41", x"56", x"C5", x"44", x"45", x"C6",
x"50", x"4F", x"4B", x"C5", x"50", x"52", x"49", x"4E",
x"D4", x"43", x"4F", x"4E", x"D4", x"4C", x"49", x"53",
x"D4", x"43", x"4C", x"45", x"41", x"D2", x"4E", x"45",
x"D7", x"54", x"41", x"42", x"A8", x"54", x"CF", x"46",
x"CE", x"53", x"50", x"43", x"A8", x"54", x"48", x"45",
x"CE", x"4E", x"4F", x"D4", x"53", x"54", x"45", x"D0",
x"AB", x"AD", x"AA", x"AF", x"E0", x"41", x"4E", x"C4",
x"4F", x"D2", x"BE", x"BD", x"BC", x"53", x"47", x"CE",
x"49", x"4E", x"D4", x"41", x"42", x"D3", x"55", x"53",
x"D2", x"46", x"52", x"C5", x"50", x"4F", x"D3", x"53",
x"51", x"D2", x"52", x"4E", x"C4", x"4C", x"4F", x"C7",
x"45", x"58", x"D0", x"43", x"4F", x"D3", x"53", x"49",
x"CE", x"54", x"41", x"CE", x"41", x"54", x"CE", x"50",
x"45", x"45", x"CB", x"4C", x"45", x"CE", x"53", x"54",
x"52", x"A4", x"56", x"41", x"CC", x"41", x"53", x"C3",
x"43", x"48", x"52", x"A4", x"4C", x"45", x"46", x"54",
x"A4", x"52", x"49", x"47", x"48", x"54", x"A4", x"4D",
x"49", x"44", x"A4", x"00", x"4E", x"46", x"53", x"4E",
x"52", x"47", x"4E", x"50", x"46", x"50", x"52", x"4F",
x"4D", x"50", x"4E", x"4E", x"50", x"50", x"44", x"44",
x"2F", x"30", x"50", x"4E", x"50", x"54", x"44", x"4E",
x"49", x"4B", x"4E", x"44", x"44", x"46", x"20", x"47",
x"52", x"45", x"5E", x"4B", x"41", x"00", x"20", x"55",
x"20", x"00", x"0D", x"0A", x"3E", x"0D", x"0A", x"00",
x"00", x"0D", x"0A", x"20", x"53", x"54", x"4F", x"50",
x"00", x"BA", x"E8", x"E8", x"E8", x"E8", x"BD", x"01",
x"01", x"C9", x"81", x"D0", x"21", x"A5", x"98", x"D0",
x"0A", x"BD", x"02", x"01", x"85", x"97", x"BD", x"03",
x"01", x"85", x"98", x"DD", x"03", x"01", x"D0", x"07",
x"A5", x"97", x"DD", x"02", x"01", x"F0", x"07", x"8A",
x"18", x"69", x"10", x"AA", x"D0", x"D8", x"60", x"20",
x"1F", x"C2", x"85", x"7F", x"84", x"80", x"38", x"A5",
x"A6", x"E5", x"AA", x"85", x"71", x"A8", x"A5", x"A7",
x"E5", x"AB", x"AA", x"E8", x"98", x"F0", x"23", x"A5",
x"A6", x"38", x"E5", x"71", x"85", x"A6", x"B0", x"03",
x"C6", x"A7", x"38", x"A5", x"A4", x"E5", x"71", x"85",
x"A4", x"B0", x"08", x"C6", x"A5", x"90", x"04", x"B1",
x"A6", x"91", x"A4", x"88", x"D0", x"F9", x"B1", x"A6",
x"91", x"A4", x"C6", x"A7", x"C6", x"A5", x"CA", x"D0",
x"F2", x"60", x"0A", x"69", x"33", x"B0", x"35", x"85",
x"71", x"BA", x"E4", x"71", x"90", x"2E", x"60", x"C4",
x"82", x"90", x"28", x"D0", x"04", x"C5", x"81", x"90",
x"22", x"48", x"A2", x"08", x"98", x"48", x"B5", x"A3",
x"CA", x"10", x"FA", x"20", x"47", x"D1", x"A2", x"F8",
x"68", x"95", x"AC", x"E8", x"30", x"FA", x"68", x"A8",
x"68", x"C4", x"82", x"90", x"06", x"D0", x"05", x"C5",
x"81", x"58", x"01", x"60", x"A2", x"0C", x"46", x"64",
x"20", x"6C", x"C8", x"20", x"E3", x"C8", x"BD", x"64",
x"C1", x"20", x"E5", x"C8", x"BD", x"65", x"C1", x"20",
x"E5", x"C8", x"20", x"91", x"C4", x"A9", x"86", x"A0",
x"C1", x"20", x"C3", x"C8", x"A4", x"88", x"C8", x"F0",
x"03", x"20", x"53", x"D9", x"46", x"64", x"A9", x"92",
x"A0", x"C1", x"20", x"03", x"00", x"20", x"57", x"C3",
x"86", x"C3", x"84", x"C4", x"20", x"BC", x"00", x"F0",
x"F4", x"A2", x"FF", x"86", x"88", x"90", x"06", x"20",
x"A6", x"C3", x"4C", x"F6", x"C5", x"20", x"7F", x"C7",
x"20", x"A6", x"C3", x"84", x"5D", x"20", x"32", x"C4",
x"90", x"44", x"A0", x"01", x"B1", x"AA", x"85", x"72",
x"A5", x"7B", x"85", x"71", x"A5", x"AB", x"85", x"74",
x"A5", x"AA", x"88", x"F1", x"AA", x"18", x"65", x"7B",
x"85", x"7B", x"85", x"73", x"A5", x"7C", x"69", x"FF",
x"85", x"7C", x"E5", x"AB", x"AA", x"38", x"A5", x"AA",
x"E5", x"7B", x"A8", x"B0", x"03", x"E8", x"C6", x"74",
x"18", x"65", x"71", x"90", x"03", x"C6", x"72", x"18",
x"B1", x"71", x"91", x"73", x"C8", x"D0", x"F9", x"E6",
x"72", x"E6", x"74", x"CA", x"D0", x"F2", x"A5", x"13",
x"F0", x"2F", x"A5", x"85", x"A4", x"86", x"85", x"81",
x"84", x"82", x"A5", x"7B", x"85", x"A6", x"65", x"5D",
x"85", x"A4", x"A4", x"7C", x"84", x"A7", x"90", x"01",
x"C8", x"84", x"A5", x"20", x"CF", x"C1", x"A5", x"7F",
x"A4", x"80", x"85", x"7B", x"84", x"7C", x"A4", x"5D",
x"88", x"B9", x"0F", x"00", x"91", x"AA", x"88", x"10",
x"F8", x"20", x"77", x"C4", x"A5", x"79", x"A4", x"7A",
x"85", x"71", x"84", x"72", x"18", x"A0", x"01", x"B1",
x"71", x"D0", x"03", x"4C", x"7D", x"C2", x"A0", x"04",
x"C8", x"B1", x"71", x"D0", x"FB", x"C8", x"98", x"65",
x"71", x"AA", x"A0", x"00", x"91", x"71", x"A5", x"72",
x"69", x"00", x"C8", x"91", x"71", x"86", x"71", x"85",
x"72", x"90", x"DA", x"20", x"E5", x"C8", x"CA", x"10",
x"08", x"20", x"E5", x"C8", x"20", x"6C", x"C8", x"A2",
x"00", x"20", x"86", x"C3", x"C9", x"0D", x"F0", x"23",
x"C9", x"40", x"F0", x"F0", x"C9", x"08", x"D0", x"05",
x"CA", x"30", x"0E", x"C6", x"0E", x"C9", x"20", x"90",
x"E8", x"E6", x"0E", x"E0", x"47", x"B0", x"05", x"95",
x"13", x"E8", x"D0", x"DD", x"A9", x"07", x"20", x"E5",
x"C8", x"D0", x"D6", x"4C", x"66", x"C8", x"20", x"EE",
x"FF", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"29",
x"FF", x"C9", x"1E", x"D0", x"08", x"48", x"A5", x"64",
x"49", x"FF", x"85", x"64", x"68", x"60", x"A6", x"C3",
x"A0", x"04", x"84", x"60", x"B5", x"00", x"C9", x"20",
x"F0", x"3A", x"85", x"5C", x"C9", x"22", x"F0", x"58",
x"24", x"60", x"70", x"30", x"C9", x"3F", x"D0", x"04",
x"A9", x"97", x"D0", x"28", x"C9", x"30", x"90", x"04",
x"C9", x"3C", x"90", x"20", x"84", x"BA", x"A0", x"00",
x"84", x"5D", x"88", x"86", x"C3", x"CA", x"C8", x"E8",
x"B5", x"00", x"C9", x"20", x"F0", x"F9", x"38", x"F9",
x"84", x"C0", x"F0", x"F2", x"C9", x"80", x"D0", x"2F",
x"05", x"5D", x"A4", x"BA", x"E8", x"C8", x"99", x"0E",
x"00", x"B9", x"0E", x"00", x"F0", x"34", x"38", x"E9",
x"3A", x"F0", x"04", x"C9", x"49", x"D0", x"02", x"85",
x"60", x"38", x"E9", x"54", x"D0", x"A6", x"85", x"5C",
x"B5", x"00", x"F0", x"E0", x"C5", x"5C", x"F0", x"DC",
x"C8", x"99", x"0E", x"00", x"E8", x"D0", x"F1", x"A6",
x"C3", x"E6", x"5D", x"C8", x"B9", x"83", x"C0", x"10",
x"FA", x"B9", x"84", x"C0", x"D0", x"B2", x"B5", x"00",
x"10", x"C0", x"99", x"10", x"00", x"A9", x"12", x"85",
x"C3", x"60", x"A5", x"79", x"A6", x"7A", x"A0", x"01",
x"85", x"AA", x"86", x"AB", x"B1", x"AA", x"F0", x"1F",
x"C8", x"C8", x"A5", x"12", x"D1", x"AA", x"90", x"18",
x"F0", x"03", x"88", x"D0", x"09", x"A5", x"11", x"88",
x"D1", x"AA", x"90", x"0C", x"F0", x"0A", x"88", x"B1",
x"AA", x"AA", x"88", x"B1", x"AA", x"B0", x"D7", x"18",
x"60", x"D0", x"FD", x"A9", x"00", x"A8", x"91", x"79",
x"C8", x"91", x"79", x"A5", x"79", x"69", x"02", x"85",
x"7B", x"A5", x"7A", x"69", x"00", x"85", x"7C", x"20",
x"A7", x"C4", x"A5", x"85", x"A4", x"86", x"85", x"81",
x"84", x"82", x"A5", x"7B", x"A4", x"7C", x"85", x"7D",
x"84", x"7E", x"85", x"7F", x"84", x"80", x"20", x"1A",
x"C6", x"A2", x"68", x"86", x"65", x"68", x"8D", x"FD",
x"01", x"68", x"8D", x"FE", x"01", x"A2", x"FC", x"9A",
x"A9", x"00", x"85", x"8C", x"85", x"61", x"60", x"18",
x"A5", x"79", x"69", x"FF", x"85", x"C3", x"A5", x"7A",
x"69", x"FF", x"85", x"C4", x"60", x"90", x"06", x"F0",
x"04", x"C9", x"A4", x"D0", x"F7", x"20", x"7F", x"C7",
x"20", x"32", x"C4", x"20", x"C2", x"00", x"F0", x"0C",
x"C9", x"A4", x"D0", x"94", x"20", x"BC", x"00", x"20",
x"7F", x"C7", x"D0", x"8C", x"68", x"68", x"A5", x"11",
x"05", x"12", x"D0", x"06", x"A9", x"FF", x"85", x"11",
x"85", x"12", x"A0", x"01", x"84", x"60", x"B1", x"AA",
x"F0", x"41", x"20", x"29", x"C6", x"20", x"6C", x"C8",
x"C8", x"B1", x"AA", x"AA", x"C8", x"B1", x"AA", x"C5",
x"12", x"D0", x"04", x"E4", x"11", x"F0", x"02", x"B0",
x"2A", x"84", x"97", x"20", x"5E", x"D9", x"A9", x"20",
x"A4", x"97", x"29", x"7F", x"20", x"E5", x"C8", x"C9",
x"22", x"D0", x"06", x"A5", x"60", x"49", x"FF", x"85",
x"60", x"C8", x"B1", x"AA", x"D0", x"10", x"A8", x"B1",
x"AA", x"AA", x"C8", x"B1", x"AA", x"86", x"AA", x"85",
x"AB", x"D0", x"B7", x"4C", x"74", x"C2", x"10", x"DC",
x"C9", x"FF", x"F0", x"D8", x"24", x"60", x"30", x"D4",
x"38", x"E9", x"7F", x"AA", x"84", x"97", x"A0", x"FF",
x"CA", x"F0", x"08", x"C8", x"B9", x"84", x"C0", x"10",
x"FA", x"30", x"F5", x"C8", x"B9", x"84", x"C0", x"30",
x"B7", x"20", x"E5", x"C8", x"D0", x"F5", x"A9", x"80",
x"85", x"61", x"20", x"B9", x"C7", x"20", x"A1", x"C1",
x"D0", x"05", x"8A", x"69", x"0D", x"AA", x"9A", x"68",
x"68", x"A9", x"08", x"20", x"12", x"C2", x"20", x"1A",
x"C7", x"18", x"98", x"65", x"C3", x"48", x"A5", x"C4",
x"69", x"00", x"48", x"A5", x"88", x"48", x"A5", x"87",
x"48", x"A9", x"9D", x"20", x"03", x"CC", x"20", x"B0",
x"CA", x"20", x"AD", x"CA", x"A5", x"B0", x"09", x"7F",
x"25", x"AD", x"85", x"AD", x"A9", x"9F", x"A0", x"C5",
x"85", x"71", x"84", x"72", x"4C", x"66", x"CB", x"A9",
x"9C", x"A0", x"D5", x"20", x"4B", x"D7", x"20", x"C2",
x"00", x"C9", x"A2", x"D0", x"06", x"20", x"BC", x"00",
x"20", x"AD", x"CA", x"20", x"CA", x"D7", x"20", x"5B",
x"CB", x"A5", x"98", x"48", x"A5", x"97", x"48", x"A9",
x"81", x"48", x"20", x"29", x"C6", x"A5", x"C3", x"A4",
x"C4", x"F0", x"06", x"85", x"8B", x"84", x"8C", x"A0",
x"00", x"B1", x"C3", x"F0", x"07", x"C9", x"3A", x"F0",
x"1D", x"4C", x"0C", x"CC", x"A0", x"02", x"B1", x"C3",
x"18", x"F0", x"6E", x"C8", x"B1", x"C3", x"85", x"87",
x"C8", x"B1", x"C3", x"85", x"88", x"98", x"65", x"C3",
x"85", x"C3", x"90", x"02", x"E6", x"C4", x"20", x"BC",
x"00", x"20", x"FF", x"C5", x"4C", x"C2", x"C5", x"F0",
x"79", x"38", x"E9", x"80", x"B0", x"03", x"4C", x"B9",
x"C7", x"C9", x"1C", x"B0", x"CC", x"0A", x"A8", x"B9",
x"01", x"C0", x"48", x"B9", x"00", x"C0", x"48", x"4C",
x"BC", x"00", x"38", x"A5", x"79", x"E9", x"01", x"A4",
x"7A", x"B0", x"01", x"88", x"85", x"8F", x"84", x"90",
x"60", x"2C", x"11", x"02", x"10", x"FA", x"20", x"0F",
x"E6", x"F0", x"F5", x"20", x"86", x"C3", x"C9", x"03",
x"B0", x"01", x"18", x"D0", x"3D", x"A5", x"C3", x"A4",
x"C4", x"F0", x"0C", x"85", x"8B", x"84", x"8C", x"A5",
x"87", x"A4", x"88", x"85", x"89", x"84", x"8A", x"68",
x"68", x"A9", x"99", x"A0", x"C1", x"A2", x"00", x"86",
x"64", x"90", x"03", x"4C", x"69", x"C2", x"4C", x"74",
x"C2", x"D0", x"17", x"A2", x"1E", x"A4", x"8C", x"D0",
x"03", x"4C", x"4E", x"C2", x"A5", x"8B", x"85", x"C3",
x"84", x"C4", x"A5", x"89", x"A4", x"8A", x"85", x"87",
x"84", x"88", x"60", x"20", x"AE", x"D3", x"D0", x"FA",
x"E8", x"E0", x"0A", x"B0", x"04", x"CA", x"86", x"0D",
x"60", x"4C", x"88", x"CE", x"D0", x"EC", x"4C", x"7A",
x"C4", x"D0", x"03", x"4C", x"77", x"C4", x"20", x"7A",
x"C4", x"4C", x"B0", x"C6", x"A9", x"03", x"20", x"12",
x"C2", x"A5", x"C4", x"48", x"A5", x"C3", x"48", x"A5",
x"88", x"48", x"A5", x"87", x"48", x"A9", x"8C", x"48",
x"20", x"C2", x"00", x"20", x"B9", x"C6", x"4C", x"C2",
x"C5", x"20", x"7F", x"C7", x"20", x"1D", x"C7", x"A5",
x"88", x"C5", x"12", x"B0", x"0B", x"98", x"38", x"65",
x"C3", x"A6", x"C4", x"90", x"07", x"E8", x"B0", x"04",
x"A5", x"79", x"A6", x"7A", x"20", x"36", x"C4", x"90",
x"1E", x"A5", x"AA", x"E9", x"01", x"85", x"C3", x"A5",
x"AB", x"E9", x"00", x"85", x"C4", x"60", x"D0", x"FD",
x"A9", x"FF", x"85", x"97", x"20", x"A1", x"C1", x"9A",
x"C9", x"8C", x"F0", x"0B", x"A2", x"04", x"2C", x"A2",
x"0E", x"4C", x"4E", x"C2", x"4C", x"0C", x"CC", x"68",
x"68", x"85", x"87", x"68", x"85", x"88", x"68", x"85",
x"C3", x"68", x"85", x"C4", x"20", x"1A", x"C7", x"98",
x"18", x"65", x"C3", x"85", x"C3", x"90", x"02", x"E6",
x"C4", x"60", x"A2", x"3A", x"2C", x"A2", x"00", x"86",
x"5B", x"A0", x"00", x"84", x"5C", x"A5", x"5C", x"A6",
x"5B", x"85", x"5B", x"86", x"5C", x"B1", x"C3", x"F0",
x"E8", x"C5", x"5C", x"F0", x"E4", x"C8", x"C9", x"22",
x"F0", x"EB", x"D0", x"F1", x"20", x"C1", x"CA", x"20",
x"C2", x"00", x"C9", x"88", x"F0", x"05", x"A9", x"A0",
x"20", x"03", x"CC", x"A5", x"AC", x"D0", x"05", x"20",
x"1D", x"C7", x"F0", x"BB", x"20", x"C2", x"00", x"B0",
x"03", x"4C", x"B9", x"C6", x"4C", x"FF", x"C5", x"20",
x"AE", x"D3", x"48", x"C9", x"8C", x"F0", x"04", x"C9",
x"88", x"D0", x"91", x"C6", x"AF", x"D0", x"04", x"68",
x"4C", x"02", x"C6", x"20", x"BC", x"00", x"20", x"7F",
x"C7", x"C9", x"2C", x"F0", x"EE", x"68", x"60", x"A2",
x"00", x"86", x"11", x"86", x"12", x"B0", x"F7", x"E9",
x"2F", x"85", x"5B", x"A5", x"12", x"85", x"71", x"C9",
x"19", x"B0", x"D4", x"A5", x"11", x"0A", x"26", x"71",
x"0A", x"26", x"71", x"65", x"11", x"85", x"11", x"A5",
x"71", x"65", x"12", x"85", x"12", x"06", x"11", x"26",
x"12", x"A5", x"11", x"65", x"5B", x"85", x"11", x"90",
x"02", x"E6", x"12", x"20", x"BC", x"00", x"4C", x"85",
x"C7", x"20", x"0B", x"CD", x"85", x"97", x"84", x"98",
x"A9", x"AB", x"20", x"03", x"CC", x"A5", x"5F", x"48",
x"20", x"C1", x"CA", x"68", x"2A", x"20", x"B3", x"CA",
x"D0", x"03", x"4C", x"74", x"D7", x"A0", x"02", x"B1",
x"AE", x"C5", x"82", x"90", x"17", x"D0", x"07", x"88",
x"B1", x"AE", x"C5", x"81", x"90", x"0E", x"A4", x"AF",
x"C4", x"7C", x"90", x"08", x"D0", x"0D", x"A5", x"AE",
x"C5", x"7B", x"B0", x"07", x"A5", x"AE", x"A4", x"AF",
x"4C", x"11", x"C8", x"A0", x"00", x"B1", x"AE", x"20",
x"9C", x"D0", x"A5", x"9E", x"A4", x"9F", x"85", x"B8",
x"84", x"B9", x"20", x"8A", x"D2", x"A9", x"AC", x"A0",
x"00", x"85", x"9E", x"84", x"9F", x"20", x"EB", x"D2",
x"A0", x"00", x"B1", x"9E", x"91", x"97", x"C8", x"B1",
x"9E", x"91", x"97", x"C8", x"B1", x"9E", x"91", x"97",
x"60", x"20", x"C6", x"C8", x"20", x"C2", x"00", x"F0",
x"3B", x"F0", x"57", x"C9", x"9C", x"F0", x"6B", x"C9",
x"9F", x"F0", x"67", x"C9", x"2C", x"F0", x"4C", x"C9",
x"3B", x"F0", x"7A", x"20", x"C1", x"CA", x"24", x"5F",
x"30", x"DF", x"20", x"6E", x"D9", x"20", x"AE", x"D0",
x"A0", x"00", x"B1", x"AE", x"18", x"65", x"0E", x"C5",
x"0F", x"90", x"03", x"20", x"6C", x"C8", x"20", x"C6",
x"C8", x"20", x"E0", x"C8", x"D0", x"C6", x"A0", x"00",
x"94", x"13", x"A2", x"12", x"A9", x"0D", x"85", x"0E",
x"20", x"E5", x"C8", x"A9", x"0A", x"20", x"E5", x"C8",
x"8A", x"48", x"A6", x"0D", x"F0", x"08", x"A9", x"00",
x"20", x"E5", x"C8", x"CA", x"D0", x"FA", x"86", x"0E",
x"68", x"AA", x"60", x"A5", x"0E", x"C5", x"10", x"90",
x"06", x"20", x"6C", x"C8", x"4C", x"BD", x"C8", x"38",
x"E9", x"0E", x"B0", x"FC", x"49", x"FF", x"69", x"01",
x"D0", x"14", x"48", x"20", x"AB", x"D3", x"C9", x"29",
x"D0", x"66", x"68", x"C9", x"9C", x"D0", x"08", x"8A",
x"E5", x"0E", x"90", x"09", x"F0", x"07", x"AA", x"20",
x"E0", x"C8", x"CA", x"D0", x"FA", x"20", x"BC", x"00",
x"4C", x"31", x"C8", x"20", x"AE", x"D0", x"20", x"B6",
x"D2", x"AA", x"A0", x"00", x"E8", x"CA", x"F0", x"BA",
x"B1", x"71", x"20", x"E5", x"C8", x"C8", x"C9", x"0D",
x"D0", x"F3", x"20", x"78", x"C8", x"4C", x"CD", x"C8",
x"A9", x"20", x"2C", x"A9", x"3F", x"24", x"64", x"30",
x"18", x"48", x"C9", x"20", x"90", x"0B", x"A5", x"0E",
x"C5", x"0F", x"D0", x"03", x"20", x"6C", x"C8", x"E6",
x"0E", x"68", x"20", x"F1", x"FF", x"EA", x"EA", x"EA",
x"EA", x"29", x"FF", x"60", x"A5", x"62", x"F0", x"0B",
x"A5", x"8D", x"A4", x"8E", x"85", x"87", x"84", x"88",
x"4C", x"0C", x"CC", x"A9", x"2D", x"A0", x"CA", x"20",
x"C3", x"C8", x"A5", x"8B", x"A4", x"8C", x"85", x"C3",
x"84", x"C4", x"60", x"46", x"64", x"C9", x"22", x"D0",
x"0B", x"20", x"C1", x"CB", x"A9", x"3B", x"20", x"03",
x"CC", x"20", x"C6", x"C8", x"20", x"D4", x"CF", x"A9",
x"2C", x"85", x"12", x"20", x"46", x"C9", x"A5", x"13",
x"D0", x"12", x"18", x"4C", x"47", x"C6", x"20", x"E3",
x"C8", x"20", x"E0", x"C8", x"4C", x"57", x"C3", x"A6",
x"8F", x"A4", x"90", x"A9", x"98", x"85", x"62", x"86",
x"91", x"84", x"92", x"20", x"0B", x"CD", x"85", x"97",
x"84", x"98", x"A5", x"C3", x"A4", x"C4", x"85", x"11",
x"84", x"12", x"A6", x"91", x"A4", x"92", x"86", x"C3",
x"84", x"C4", x"20", x"C2", x"00", x"D0", x"0E", x"24",
x"62", x"30", x"62", x"20", x"E3", x"C8", x"20", x"46",
x"C9", x"86", x"C3", x"84", x"C4", x"20", x"BC", x"00",
x"24", x"5F", x"10", x"24", x"85", x"5B", x"C9", x"22",
x"F0", x"07", x"A9", x"3A", x"85", x"5B", x"A9", x"2C",
x"18", x"85", x"5C", x"A5", x"C3", x"A4", x"C4", x"69",
x"00", x"90", x"01", x"C8", x"20", x"B4", x"D0", x"20",
x"F3", x"D3", x"20", x"D5", x"C7", x"4C", x"B6", x"C9",
x"20", x"87", x"D8", x"20", x"74", x"D7", x"20", x"C2",
x"00", x"F0", x"07", x"C9", x"2C", x"F0", x"03", x"4C",
x"04", x"C9", x"A5", x"C3", x"A4", x"C4", x"85", x"91",
x"84", x"92", x"A5", x"11", x"A4", x"12", x"85", x"C3",
x"84", x"C4", x"20", x"C2", x"00", x"F0", x"2C", x"20",
x"01", x"CC", x"4C", x"5B", x"C9", x"20", x"1A", x"C7",
x"C8", x"AA", x"D0", x"12", x"A2", x"06", x"C8", x"B1",
x"C3", x"F0", x"69", x"C8", x"B1", x"C3", x"85", x"8D",
x"C8", x"B1", x"C3", x"C8", x"85", x"8E", x"B1", x"C3",
x"AA", x"20", x"0F", x"C7", x"E0", x"83", x"D0", x"DD",
x"4C", x"85", x"C9", x"A5", x"91", x"A4", x"92", x"A6",
x"62", x"F0", x"03", x"4C", x"24", x"C6", x"A0", x"00",
x"B1", x"91", x"F0", x"07", x"A9", x"1C", x"A0", x"CA",
x"4C", x"C3", x"C8", x"60", x"3F", x"50", x"52", x"45",
x"56", x"49", x"5E", x"45", x"20", x"55", x"4C", x"41",
x"5A", x"41", x"0D", x"0A", x"00", x"20", x"3F", x"20",
x"50", x"4F", x"4E", x"4F", x"56", x"49", x"20", x"55",
x"50", x"49", x"53", x"20", x"20", x"0D", x"0A", x"00",
x"D0", x"04", x"A0", x"00", x"F0", x"03", x"20", x"0B",
x"CD", x"85", x"97", x"84", x"98", x"20", x"A1", x"C1",
x"F0", x"04", x"A2", x"00", x"F0", x"68", x"9A", x"E8",
x"E8", x"E8", x"E8", x"8A", x"E8", x"E8", x"E8", x"E8",
x"E8", x"86", x"73", x"A0", x"01", x"20", x"4B", x"D7",
x"BA", x"BD", x"08", x"01", x"85", x"B0", x"A5", x"97",
x"A4", x"98", x"20", x"6C", x"D4", x"20", x"74", x"D7",
x"A0", x"01", x"20", x"FA", x"D7", x"BA", x"38", x"FD",
x"08", x"01", x"F0", x"17", x"BD", x"0D", x"01", x"85",
x"87", x"BD", x"0E", x"01", x"85", x"88", x"BD", x"10",
x"01", x"85", x"C3", x"BD", x"0F", x"01", x"85", x"C4",
x"4C", x"C2", x"C5", x"8A", x"69", x"0F", x"AA", x"9A",
x"20", x"C2", x"00", x"C9", x"2C", x"D0", x"F1", x"20",
x"BC", x"00", x"20", x"46", x"CA", x"20", x"C1", x"CA",
x"18", x"24", x"38", x"24", x"5F", x"30", x"03", x"B0",
x"03", x"60", x"B0", x"FD", x"A2", x"18", x"4C", x"4E",
x"C2", x"A6", x"C3", x"D0", x"02", x"C6", x"C4", x"C6",
x"C3", x"A2", x"00", x"24", x"48", x"8A", x"48", x"A9",
x"01", x"20", x"12", x"C2", x"20", x"A0", x"CB", x"A9",
x"00", x"85", x"9B", x"20", x"C2", x"00", x"38", x"E9",
x"AA", x"90", x"17", x"C9", x"03", x"B0", x"13", x"C9",
x"01", x"2A", x"49", x"01", x"45", x"9B", x"C5", x"9B",
x"90", x"61", x"85", x"9B", x"20", x"BC", x"00", x"4C",
x"DE", x"CA", x"A6", x"9B", x"D0", x"2C", x"B0", x"78",
x"69", x"07", x"90", x"74", x"65", x"5F", x"D0", x"03",
x"4C", x"4D", x"D2", x"69", x"FF", x"85", x"71", x"0A",
x"65", x"71", x"A8", x"68", x"D9", x"66", x"C0", x"B0",
x"64", x"20", x"B0", x"CA", x"48", x"20", x"43", x"CB",
x"68", x"A4", x"99", x"10", x"17", x"AA", x"F0", x"53",
x"D0", x"5C", x"46", x"5F", x"8A", x"2A", x"A6", x"C3",
x"D0", x"02", x"C6", x"C4", x"C6", x"C3", x"A0", x"1B",
x"85", x"9B", x"D0", x"D7", x"D9", x"66", x"C0", x"B0",
x"45", x"90", x"D9", x"B9", x"68", x"C0", x"48", x"B9",
x"67", x"C0", x"48", x"20", x"56", x"CB", x"A5", x"9B",
x"4C", x"CC", x"CA", x"4C", x"0C", x"CC", x"A5", x"B0",
x"BE", x"66", x"C0", x"A8", x"68", x"85", x"71", x"E6",
x"71", x"68", x"85", x"72", x"98", x"48", x"20", x"BA",
x"D7", x"A5", x"AF", x"48", x"A5", x"AE", x"48", x"A5",
x"AD", x"48", x"A5", x"AC", x"48", x"6C", x"71", x"00",
x"A0", x"FF", x"68", x"F0", x"20", x"C9", x"64", x"F0",
x"03", x"20", x"B0", x"CA", x"84", x"99", x"68", x"4A",
x"85", x"63", x"68", x"85", x"B3", x"68", x"85", x"B4",
x"68", x"85", x"B5", x"68", x"85", x"B6", x"68", x"85",
x"B7", x"45", x"B0", x"85", x"B8", x"A5", x"AC", x"60",
x"A9", x"00", x"85", x"5F", x"20", x"BC", x"00", x"B0",
x"03", x"4C", x"87", x"D8", x"20", x"81", x"CD", x"B0",
x"67", x"C9", x"2E", x"F0", x"F4", x"C9", x"A4", x"F0",
x"58", x"C9", x"A3", x"F0", x"E7", x"C9", x"22", x"D0",
x"0F", x"A5", x"C3", x"A4", x"C4", x"69", x"00", x"90",
x"01", x"C8", x"20", x"AE", x"D0", x"4C", x"F3", x"D3",
x"C9", x"A1", x"D0", x"13", x"A0", x"18", x"D0", x"3B",
x"20", x"05", x"CE", x"A5", x"AF", x"49", x"FF", x"A8",
x"A5", x"AE", x"49", x"FF", x"4C", x"C1", x"CF", x"C9",
x"9E", x"D0", x"03", x"4C", x"1E", x"D0", x"C9", x"AD",
x"90", x"03", x"4C", x"27", x"CC", x"20", x"FE", x"CB",
x"20", x"C1", x"CA", x"A9", x"29", x"2C", x"A9", x"28",
x"2C", x"A9", x"2C", x"A0", x"00", x"D1", x"C3", x"D0",
x"03", x"4C", x"BC", x"00", x"A2", x"02", x"4C", x"4E",
x"C2", x"A0", x"15", x"68", x"68", x"4C", x"1D", x"CB",
x"20", x"0B", x"CD", x"85", x"AE", x"84", x"AF", x"A6",
x"5F", x"F0", x"01", x"60", x"4C", x"4B", x"D7", x"0A",
x"48", x"AA", x"20", x"BC", x"00", x"E0", x"81", x"90",
x"20", x"20", x"FE", x"CB", x"20", x"C1", x"CA", x"20",
x"01", x"CC", x"20", x"B2", x"CA", x"68", x"AA", x"A5",
x"AF", x"48", x"A5", x"AE", x"48", x"8A", x"48", x"20",
x"AE", x"D3", x"68", x"A8", x"8A", x"48", x"4C", x"56",
x"CC", x"20", x"F5", x"CB", x"68", x"A8", x"B9", x"DE",
x"BF", x"85", x"A2", x"B9", x"DF", x"BF", x"85", x"A3",
x"20", x"A1", x"00", x"4C", x"B0", x"CA", x"A0", x"FF",
x"2C", x"A0", x"00", x"84", x"5D", x"20", x"05", x"CE",
x"A5", x"AE", x"45", x"5D", x"85", x"5B", x"A5", x"AF",
x"45", x"5D", x"85", x"5C", x"20", x"9B", x"D7", x"20",
x"05", x"CE", x"A5", x"AF", x"45", x"5D", x"25", x"5C",
x"45", x"5D", x"A8", x"A5", x"AE", x"45", x"5D", x"25",
x"5B", x"45", x"5D", x"4C", x"C1", x"CF", x"20", x"B3",
x"CA", x"B0", x"13", x"A5", x"B7", x"09", x"7F", x"25",
x"B4", x"85", x"B4", x"A9", x"B3", x"A0", x"00", x"20",
x"F8", x"D7", x"AA", x"4C", x"E1", x"CC", x"A9", x"00",
x"85", x"5F", x"C6", x"9B", x"20", x"B6", x"D2", x"85",
x"AC", x"86", x"AD", x"84", x"AE", x"A5", x"B5", x"A4",
x"B6", x"20", x"BA", x"D2", x"86", x"B5", x"84", x"B6",
x"AA", x"38", x"E5", x"AC", x"F0", x"08", x"A9", x"01",
x"90", x"04", x"A6", x"AC", x"A9", x"FF", x"85", x"B0",
x"A0", x"FF", x"E8", x"C8", x"CA", x"D0", x"07", x"A6",
x"B0", x"30", x"0F", x"18", x"90", x"0C", x"B1", x"B5",
x"D1", x"AD", x"F0", x"EF", x"A2", x"FF", x"B0", x"02",
x"A2", x"01", x"E8", x"8A", x"2A", x"25", x"63", x"F0",
x"02", x"A9", x"FF", x"4C", x"DB", x"D7", x"20", x"01",
x"CC", x"AA", x"20", x"10", x"CD", x"20", x"C2", x"00",
x"D0", x"F4", x"60", x"A2", x"00", x"20", x"C2", x"00",
x"86", x"5E", x"85", x"93", x"20", x"C2", x"00", x"20",
x"81", x"CD", x"B0", x"03", x"4C", x"0C", x"CC", x"A2",
x"00", x"86", x"5F", x"20", x"BC", x"00", x"90", x"05",
x"20", x"81", x"CD", x"90", x"0B", x"AA", x"20", x"BC",
x"00", x"90", x"FB", x"20", x"81", x"CD", x"B0", x"F6",
x"C9", x"24", x"D0", x"0B", x"A9", x"FF", x"85", x"5F",
x"8A", x"09", x"80", x"AA", x"20", x"BC", x"00", x"86",
x"94", x"38", x"05", x"61", x"E9", x"28", x"D0", x"03",
x"4C", x"17", x"CE", x"A9", x"00", x"85", x"61", x"A5",
x"7B", x"A6", x"7C", x"A0", x"00", x"86", x"AB", x"85",
x"AA", x"E4", x"7E", x"D0", x"04", x"C5", x"7D", x"F0",
x"22", x"A5", x"93", x"D1", x"AA", x"D0", x"08", x"A5",
x"94", x"C8", x"D1", x"AA", x"F0", x"61", x"88", x"18",
x"A5", x"AA", x"69", x"06", x"90", x"E1", x"E8", x"D0",
x"DC", x"C9", x"41", x"90", x"05", x"E9", x"5B", x"38",
x"E9", x"A5", x"60", x"68", x"48", x"C9", x"1A", x"D0",
x"07", x"A9", x"96", x"A0", x"CD", x"60", x"00", x"00",
x"A5", x"7D", x"A4", x"7E", x"85", x"AA", x"84", x"AB",
x"A5", x"7F", x"A4", x"80", x"85", x"A6", x"84", x"A7",
x"18", x"69", x"06", x"90", x"01", x"C8", x"85", x"A4",
x"84", x"A5", x"20", x"CF", x"C1", x"A5", x"A4", x"A4",
x"A5", x"C8", x"85", x"7D", x"84", x"7E", x"A0", x"00",
x"A5", x"93", x"91", x"AA", x"C8", x"A5", x"94", x"91",
x"AA", x"A9", x"00", x"C8", x"91", x"AA", x"C8", x"91",
x"AA", x"C8", x"91", x"AA", x"C8", x"91", x"AA", x"A5",
x"AA", x"18", x"69", x"02", x"A4", x"AB", x"90", x"01",
x"C8", x"85", x"95", x"84", x"96", x"60", x"A5", x"5D",
x"0A", x"69", x"05", x"65", x"AA", x"A4", x"AB", x"90",
x"01", x"C8", x"85", x"A4", x"84", x"A5", x"60", x"90",
x"80", x"00", x"00", x"20", x"BC", x"00", x"20", x"AD",
x"CA", x"A5", x"B0", x"30", x"0D", x"A5", x"AC", x"C9",
x"90", x"90", x"09", x"A9", x"F7", x"A0", x"CD", x"20",
x"F8", x"D7", x"D0", x"74", x"4C", x"31", x"D8", x"A5",
x"5E", x"48", x"A5", x"5F", x"48", x"A0", x"00", x"98",
x"48", x"A5", x"94", x"48", x"A5", x"93", x"48", x"20",
x"FB", x"CD", x"68", x"85", x"93", x"68", x"85", x"94",
x"68", x"A8", x"BA", x"BD", x"02", x"01", x"48", x"BD",
x"01", x"01", x"48", x"A5", x"AE", x"9D", x"02", x"01",
x"A5", x"AF", x"9D", x"01", x"01", x"C8", x"20", x"C2",
x"00", x"C9", x"2C", x"F0", x"D2", x"84", x"5D", x"20",
x"FB", x"CB", x"68", x"85", x"5F", x"68", x"85", x"5E",
x"A6", x"7D", x"A5", x"7E", x"86", x"AA", x"85", x"AB",
x"C5", x"80", x"D0", x"04", x"E4", x"7F", x"F0", x"39",
x"A0", x"00", x"B1", x"AA", x"C8", x"C5", x"93", x"D0",
x"06", x"A5", x"94", x"D1", x"AA", x"F0", x"16", x"C8",
x"B1", x"AA", x"18", x"65", x"AA", x"AA", x"C8", x"B1",
x"AA", x"65", x"AB", x"90", x"D7", x"A2", x"10", x"2C",
x"A2", x"08", x"4C", x"4E", x"C2", x"A2", x"12", x"A5",
x"5E", x"D0", x"F7", x"20", x"E6", x"CD", x"A5", x"5D",
x"A0", x"04", x"D1", x"AA", x"D0", x"E7", x"4C", x"24",
x"CF", x"20", x"E6", x"CD", x"20", x"1F", x"C2", x"A9",
x"00", x"A8", x"85", x"BB", x"A2", x"04", x"86", x"BA",
x"A5", x"93", x"91", x"AA", x"C8", x"A5", x"94", x"91",
x"AA", x"A5", x"5D", x"C8", x"C8", x"C8", x"91", x"AA",
x"A2", x"0B", x"A9", x"00", x"24", x"5E", x"50", x"08",
x"68", x"18", x"69", x"01", x"AA", x"68", x"69", x"00",
x"C8", x"91", x"AA", x"C8", x"8A", x"91", x"AA", x"20",
x"7C", x"CF", x"86", x"BA", x"85", x"BB", x"A4", x"71",
x"C6", x"5D", x"D0", x"DC", x"65", x"A5", x"B0", x"5D",
x"85", x"A5", x"A8", x"8A", x"65", x"A4", x"90", x"03",
x"C8", x"F0", x"52", x"20", x"1F", x"C2", x"85", x"7F",
x"84", x"80", x"A9", x"00", x"E6", x"BB", x"A4", x"BA",
x"F0", x"05", x"88", x"91", x"A4", x"D0", x"FB", x"C6",
x"A5", x"C6", x"BB", x"D0", x"F5", x"E6", x"A5", x"38",
x"A5", x"7F", x"E5", x"AA", x"A0", x"02", x"91", x"AA",
x"A5", x"80", x"C8", x"E5", x"AB", x"91", x"AA", x"A5",
x"5E", x"D0", x"58", x"C8", x"B1", x"AA", x"85", x"5D",
x"A9", x"00", x"85", x"BA", x"85", x"BB", x"C8", x"68",
x"AA", x"85", x"AE", x"68", x"85", x"AF", x"D1", x"AA",
x"90", x"0E", x"D0", x"06", x"C8", x"8A", x"D1", x"AA",
x"90", x"07", x"4C", x"85", x"CE", x"4C", x"4C", x"C2",
x"C8", x"A5", x"BB", x"05", x"BA", x"18", x"F0", x"0A",
x"20", x"7C", x"CF", x"8A", x"65", x"AE", x"AA", x"98",
x"A4", x"71", x"65", x"AF", x"86", x"BA", x"C6", x"5D",
x"D0", x"CA", x"06", x"BA", x"2A", x"B0", x"DB", x"06",
x"BA", x"2A", x"B0", x"D6", x"A8", x"A5", x"BA", x"65",
x"A4", x"85", x"95", x"98", x"65", x"A5", x"85", x"96",
x"A8", x"A5", x"95", x"60", x"84", x"71", x"B1", x"AA",
x"85", x"76", x"88", x"B1", x"AA", x"85", x"77", x"A9",
x"10", x"85", x"A8", x"A2", x"00", x"A0", x"00", x"8A",
x"0A", x"AA", x"98", x"2A", x"A8", x"B0", x"AE", x"06",
x"BA", x"26", x"BB", x"90", x"0B", x"18", x"8A", x"65",
x"76", x"AA", x"98", x"65", x"77", x"A8", x"B0", x"9D",
x"C6", x"A8", x"D0", x"E3", x"60", x"A5", x"5F", x"F0",
x"03", x"20", x"B6", x"D2", x"20", x"47", x"D1", x"38",
x"A5", x"81", x"E5", x"7F", x"A8", x"A5", x"82", x"E5",
x"80", x"A2", x"00", x"86", x"5F", x"85", x"AD", x"84",
x"AE", x"A2", x"90", x"4C", x"E3", x"D7", x"A4", x"0E",
x"A9", x"00", x"F0", x"ED", x"A6", x"88", x"E8", x"D0",
x"A2", x"A2", x"16", x"4C", x"4E", x"C2", x"20", x"0B",
x"D0", x"20", x"D4", x"CF", x"20", x"FE", x"CB", x"A9",
x"80", x"85", x"61", x"20", x"0B", x"CD", x"20", x"B0",
x"CA", x"20", x"FB", x"CB", x"A9", x"AB", x"20", x"03",
x"CC", x"A5", x"96", x"48", x"A5", x"95", x"48", x"A5",
x"C4", x"48", x"A5", x"C3", x"48", x"20", x"0C", x"C7",
x"4C", x"7A", x"D0", x"A9", x"9E", x"20", x"03", x"CC",
x"09", x"80", x"85", x"61", x"20", x"12", x"CD", x"85",
x"9C", x"84", x"9D", x"4C", x"B0", x"CA", x"20", x"0B",
x"D0", x"A5", x"9D", x"48", x"A5", x"9C", x"48", x"20",
x"F5", x"CB", x"20", x"B0", x"CA", x"68", x"85", x"9C",
x"68", x"85", x"9D", x"A0", x"02", x"A2", x"20", x"B1",
x"9C", x"F0", x"A0", x"85", x"95", x"AA", x"C8", x"B1",
x"9C", x"85", x"96", x"B1", x"95", x"48", x"88", x"10",
x"FA", x"A4", x"96", x"20", x"78", x"D7", x"A5", x"C4",
x"48", x"A5", x"C3", x"48", x"B1", x"9C", x"85", x"C3",
x"C8", x"B1", x"9C", x"85", x"C4", x"A5", x"96", x"48",
x"A5", x"95", x"48", x"20", x"AD", x"CA", x"68", x"85",
x"9C", x"68", x"85", x"9D", x"20", x"C2", x"00", x"F0",
x"03", x"4C", x"0C", x"CC", x"68", x"85", x"C3", x"68",
x"85", x"C4", x"A0", x"00", x"68", x"91", x"9C", x"68",
x"C8", x"91", x"9C", x"68", x"C8", x"91", x"9C", x"68",
x"C8", x"91", x"9C", x"60", x"20", x"B0", x"CA", x"A0",
x"00", x"20", x"70", x"D9", x"68", x"68", x"A9", x"FF",
x"A0", x"00", x"F0", x"12", x"A6", x"AE", x"A4", x"AF",
x"86", x"9E", x"84", x"9F", x"20", x"15", x"D1", x"86",
x"AD", x"84", x"AE", x"85", x"AC", x"60", x"A2", x"22",
x"86", x"5B", x"86", x"5C", x"85", x"B8", x"84", x"B9",
x"85", x"AD", x"84", x"AE", x"A0", x"FF", x"C8", x"B1",
x"B8", x"F0", x"0C", x"C5", x"5B", x"F0", x"04", x"C5",
x"5C", x"D0", x"F3", x"C9", x"22", x"F0", x"01", x"18",
x"84", x"AC", x"98", x"65", x"B8", x"85", x"BA", x"A6",
x"B9", x"90", x"01", x"E8", x"86", x"BB", x"A5", x"B9",
x"D0", x"0B", x"98", x"20", x"9C", x"D0", x"A6", x"B8",
x"A4", x"B9", x"20", x"98", x"D2", x"A6", x"65", x"E0",
x"71", x"D0", x"05", x"A2", x"1C", x"4C", x"4E", x"C2",
x"A5", x"AC", x"95", x"00", x"A5", x"AD", x"95", x"01",
x"A5", x"AE", x"95", x"02", x"A0", x"00", x"86", x"AE",
x"84", x"AF", x"88", x"84", x"5F", x"86", x"66", x"E8",
x"E8", x"E8", x"86", x"65", x"60", x"46", x"60", x"48",
x"49", x"FF", x"38", x"65", x"81", x"A4", x"82", x"B0",
x"01", x"88", x"C4", x"80", x"90", x"11", x"D0", x"04",
x"C5", x"7F", x"90", x"0B", x"85", x"81", x"84", x"82",
x"85", x"83", x"84", x"84", x"AA", x"68", x"60", x"A2",
x"0C", x"A5", x"60", x"30", x"B8", x"20", x"47", x"D1",
x"A9", x"80", x"85", x"60", x"68", x"D0", x"D0", x"A6",
x"85", x"A5", x"86", x"86", x"81", x"85", x"82", x"A0",
x"00", x"84", x"9D", x"A5", x"7F", x"A6", x"80", x"85",
x"AA", x"86", x"AB", x"A9", x"68", x"A2", x"00", x"85",
x"71", x"86", x"72", x"C5", x"65", x"F0", x"05", x"20",
x"D9", x"D1", x"F0", x"F7", x"A9", x"06", x"85", x"A0",
x"A5", x"7B", x"A6", x"7C", x"85", x"71", x"86", x"72",
x"E4", x"7E", x"D0", x"04", x"C5", x"7D", x"F0", x"05",
x"20", x"D3", x"D1", x"F0", x"F3", x"85", x"A4", x"86",
x"A5", x"A9", x"03", x"85", x"A0", x"A5", x"A4", x"A6",
x"A5", x"E4", x"80", x"D0", x"07", x"C5", x"7F", x"D0",
x"03", x"4C", x"18", x"D2", x"85", x"71", x"86", x"72",
x"A0", x"01", x"B1", x"71", x"08", x"C8", x"B1", x"71",
x"65", x"A4", x"85", x"A4", x"C8", x"B1", x"71", x"65",
x"A5", x"85", x"A5", x"28", x"10", x"D7", x"C8", x"B1",
x"71", x"0A", x"69", x"05", x"65", x"71", x"85", x"71",
x"90", x"02", x"E6", x"72", x"A6", x"72", x"E4", x"A5",
x"D0", x"04", x"C5", x"A4", x"F0", x"C3", x"20", x"D9",
x"D1", x"F0", x"F3", x"C8", x"B1", x"71", x"10", x"30",
x"C8", x"B1", x"71", x"F0", x"2B", x"C8", x"B1", x"71",
x"AA", x"C8", x"B1", x"71", x"C5", x"82", x"90", x"06",
x"D0", x"1E", x"E4", x"81", x"B0", x"1A", x"C5", x"AB",
x"90", x"16", x"D0", x"04", x"E4", x"AA", x"90", x"10",
x"86", x"AA", x"85", x"AB", x"A5", x"71", x"A6", x"72",
x"85", x"9C", x"86", x"9D", x"A5", x"A0", x"85", x"A2",
x"A5", x"A0", x"18", x"65", x"71", x"85", x"71", x"90",
x"02", x"E6", x"72", x"A6", x"72", x"A0", x"00", x"60",
x"A6", x"9D", x"F0", x"F7", x"A5", x"A2", x"29", x"04",
x"4A", x"A8", x"85", x"A2", x"B1", x"9C", x"65", x"AA",
x"85", x"A6", x"A5", x"AB", x"69", x"00", x"85", x"A7",
x"A5", x"81", x"A6", x"82", x"85", x"A4", x"86", x"A5",
x"20", x"D6", x"C1", x"A4", x"A2", x"C8", x"A5", x"A4",
x"91", x"9C", x"AA", x"E6", x"A5", x"A5", x"A5", x"C8",
x"91", x"9C", x"4C", x"4B", x"D1", x"A5", x"AF", x"48",
x"A5", x"AE", x"48", x"20", x"A0", x"CB", x"20", x"B2",
x"CA", x"68", x"85", x"B8", x"68", x"85", x"B9", x"A0",
x"00", x"B1", x"B8", x"18", x"71", x"AE", x"90", x"05",
x"A2", x"1A", x"4C", x"4E", x"C2", x"20", x"9C", x"D0",
x"20", x"8A", x"D2", x"A5", x"9E", x"A4", x"9F", x"20",
x"BA", x"D2", x"20", x"9C", x"D2", x"A5", x"B8", x"A4",
x"B9", x"20", x"BA", x"D2", x"20", x"ED", x"D0", x"4C",
x"DB", x"CA", x"A0", x"00", x"B1", x"B8", x"48", x"C8",
x"B1", x"B8", x"AA", x"C8", x"B1", x"B8", x"A8", x"68",
x"86", x"71", x"84", x"72", x"A8", x"F0", x"0A", x"48",
x"88", x"B1", x"71", x"91", x"83", x"98", x"D0", x"F8",
x"68", x"18", x"65", x"83", x"85", x"83", x"90", x"02",
x"E6", x"84", x"60", x"20", x"B2", x"CA", x"A5", x"AE",
x"A4", x"AF", x"85", x"71", x"84", x"72", x"20", x"EB",
x"D2", x"08", x"A0", x"00", x"B1", x"71", x"48", x"C8",
x"B1", x"71", x"AA", x"C8", x"B1", x"71", x"A8", x"68",
x"28", x"D0", x"13", x"C4", x"82", x"D0", x"0F", x"E4",
x"81", x"D0", x"0B", x"48", x"18", x"65", x"81", x"85",
x"81", x"90", x"02", x"E6", x"82", x"68", x"86", x"71",
x"84", x"72", x"60", x"C4", x"67", x"D0", x"0C", x"C5",
x"66", x"D0", x"08", x"85", x"65", x"E9", x"03", x"85",
x"66", x"A0", x"00", x"60", x"20", x"B1", x"D3", x"8A",
x"48", x"A9", x"01", x"20", x"A4", x"D0", x"68", x"A0",
x"00", x"91", x"AD", x"68", x"68", x"4C", x"ED", x"D0",
x"20", x"6F", x"D3", x"D1", x"9E", x"98", x"90", x"04",
x"B1", x"9E", x"AA", x"98", x"48", x"8A", x"48", x"20",
x"A4", x"D0", x"A5", x"9E", x"A4", x"9F", x"20", x"BA",
x"D2", x"68", x"A8", x"68", x"18", x"65", x"71", x"85",
x"71", x"90", x"02", x"E6", x"72", x"98", x"20", x"9C",
x"D2", x"4C", x"ED", x"D0", x"20", x"6F", x"D3", x"18",
x"F1", x"9E", x"49", x"FF", x"4C", x"16", x"D3", x"A9",
x"FF", x"85", x"AF", x"20", x"C2", x"00", x"C9", x"29",
x"F0", x"06", x"20", x"01", x"CC", x"20", x"AE", x"D3",
x"20", x"6F", x"D3", x"CA", x"8A", x"48", x"18", x"A2",
x"00", x"F1", x"9E", x"B0", x"B8", x"49", x"FF", x"C5",
x"AF", x"90", x"B3", x"A5", x"AF", x"B0", x"AF", x"20",
x"FB", x"CB", x"68", x"85", x"A2", x"68", x"85", x"A3",
x"68", x"68", x"68", x"AA", x"68", x"85", x"9E", x"68",
x"85", x"9F", x"A0", x"00", x"8A", x"F0", x"21", x"E6",
x"A2", x"6C", x"A2", x"00", x"20", x"92", x"D3", x"4C",
x"D0", x"CF", x"20", x"B3", x"D2", x"A2", x"00", x"86",
x"5F", x"A8", x"60", x"20", x"92", x"D3", x"F0", x"08",
x"A0", x"00", x"B1", x"71", x"A8", x"4C", x"8F", x"D3",
x"4C", x"88", x"CE", x"20", x"BC", x"00", x"20", x"AD",
x"CA", x"20", x"01", x"CE", x"A6", x"AE", x"D0", x"F0",
x"A6", x"AF", x"4C", x"C2", x"00", x"20", x"92", x"D3",
x"D0", x"03", x"4C", x"F1", x"D4", x"A6", x"C3", x"A4",
x"C4", x"86", x"BA", x"84", x"BB", x"A6", x"71", x"86",
x"C3", x"18", x"65", x"71", x"85", x"73", x"A6", x"72",
x"86", x"C4", x"90", x"01", x"E8", x"86", x"74", x"A0",
x"00", x"B1", x"73", x"48", x"A9", x"00", x"91", x"73",
x"20", x"C2", x"00", x"20", x"87", x"D8", x"68", x"A0",
x"00", x"91", x"73", x"A6", x"BA", x"A4", x"BB", x"86",
x"C3", x"84", x"C4", x"60", x"20", x"AD", x"CA", x"20",
x"08", x"D4", x"20", x"01", x"CC", x"4C", x"AE", x"D3",
x"A5", x"B0", x"30", x"9C", x"A5", x"AC", x"C9", x"91",
x"B0", x"96", x"20", x"31", x"D8", x"A5", x"AE", x"A4",
x"AF", x"84", x"11", x"85", x"12", x"60", x"20", x"08",
x"D4", x"A0", x"00", x"B1", x"11", x"A8", x"4C", x"D0",
x"CF", x"20", x"FC", x"D3", x"8A", x"A0", x"00", x"91",
x"11", x"60", x"20", x"FC", x"D3", x"86", x"97", x"A2",
x"00", x"20", x"C2", x"00", x"F0", x"03", x"20", x"02",
x"D4", x"86", x"98", x"A0", x"00", x"B1", x"11", x"45",
x"98", x"25", x"97", x"F0", x"F8", x"60", x"A9", x"96",
x"A0", x"DA", x"4C", x"6C", x"D4", x"20", x"4D", x"D6",
x"A5", x"B0", x"49", x"FF", x"85", x"B0", x"45", x"B7",
x"85", x"B8", x"A5", x"AC", x"4C", x"6F", x"D4", x"20",
x"7B", x"D5", x"90", x"3C", x"20", x"4D", x"D6", x"D0",
x"03", x"4C", x"9B", x"D7", x"A6", x"B9", x"86", x"A3",
x"A2", x"B3", x"A5", x"B3", x"A8", x"F0", x"CE", x"38",
x"E5", x"AC", x"F0", x"24", x"90", x"12", x"84", x"AC",
x"A4", x"B7", x"84", x"B0", x"49", x"FF", x"69", x"00",
x"A0", x"00", x"84", x"A3", x"A2", x"AC", x"D0", x"04",
x"A0", x"00", x"84", x"B9", x"C9", x"F9", x"30", x"C7",
x"A8", x"A5", x"B9", x"56", x"01", x"20", x"92", x"D5",
x"24", x"B8", x"10", x"4C", x"A0", x"AC", x"E0", x"B3",
x"F0", x"02", x"A0", x"B3", x"38", x"49", x"FF", x"65",
x"A3", x"85", x"B9", x"B9", x"03", x"00", x"F5", x"03",
x"85", x"AF", x"B9", x"02", x"00", x"F5", x"02", x"85",
x"AE", x"B9", x"01", x"00", x"F5", x"01", x"85", x"AD",
x"B0", x"03", x"20", x"37", x"D5", x"A0", x"00", x"98",
x"18", x"A6", x"AD", x"D0", x"3E", x"A6", x"AE", x"86",
x"AD", x"A6", x"AF", x"86", x"AE", x"A6", x"B9", x"86",
x"AF", x"84", x"B9", x"69", x"08", x"C9", x"18", x"D0",
x"E8", x"A9", x"00", x"85", x"AC", x"85", x"B0", x"60",
x"65", x"A3", x"85", x"B9", x"A5", x"AF", x"65", x"B6",
x"85", x"AF", x"A5", x"AE", x"65", x"B5", x"85", x"AE",
x"A5", x"AD", x"65", x"B4", x"85", x"AD", x"4C", x"28",
x"D5", x"69", x"01", x"06", x"B9", x"26", x"AF", x"26",
x"AE", x"26", x"AD", x"10", x"F4", x"38", x"E5", x"AC",
x"B0", x"CF", x"49", x"FF", x"69", x"01", x"85", x"AC",
x"90", x"0C", x"E6", x"AC", x"F0", x"36", x"66", x"AD",
x"66", x"AE", x"66", x"AF", x"66", x"B9", x"60", x"A5",
x"B0", x"49", x"FF", x"85", x"B0", x"A5", x"AD", x"49",
x"FF", x"85", x"AD", x"A5", x"AE", x"49", x"FF", x"85",
x"AE", x"A5", x"AF", x"49", x"FF", x"85", x"AF", x"A5",
x"B9", x"49", x"FF", x"85", x"B9", x"E6", x"B9", x"D0",
x"0A", x"E6", x"AF", x"D0", x"06", x"E6", x"AE", x"D0",
x"02", x"E6", x"AD", x"60", x"A2", x"0A", x"4C", x"4E",
x"C2", x"A2", x"74", x"B4", x"03", x"84", x"B9", x"B4",
x"02", x"94", x"03", x"B4", x"01", x"94", x"02", x"A4",
x"B2", x"94", x"01", x"69", x"08", x"30", x"EC", x"F0",
x"EA", x"E9", x"08", x"A8", x"A5", x"B9", x"B0", x"12",
x"16", x"01", x"90", x"02", x"F6", x"01", x"76", x"01",
x"76", x"01", x"76", x"02", x"76", x"03", x"6A", x"C8",
x"D0", x"EE", x"18", x"60", x"81", x"00", x"00", x"00",
x"02", x"80", x"19", x"56", x"62", x"80", x"76", x"22",
x"F3", x"82", x"38", x"AA", x"40", x"80", x"35", x"04",
x"F3", x"81", x"35", x"04", x"F3", x"80", x"80", x"00",
x"00", x"80", x"31", x"72", x"18", x"20", x"CA", x"D7",
x"F0", x"02", x"10", x"03", x"4C", x"88", x"CE", x"A5",
x"AC", x"E9", x"7F", x"48", x"A9", x"80", x"85", x"AC",
x"A9", x"AD", x"A0", x"D5", x"20", x"6C", x"D4", x"A9",
x"B1", x"A0", x"D5", x"20", x"CA", x"D6", x"A9", x"9C",
x"A0", x"D5", x"20", x"55", x"D4", x"A9", x"A0", x"A0",
x"D5", x"20", x"6E", x"DB", x"A9", x"B5", x"A0", x"D5",
x"20", x"6C", x"D4", x"68", x"20", x"12", x"D9", x"A9",
x"B9", x"A0", x"D5", x"20", x"4D", x"D6", x"F0", x"4C",
x"20", x"73", x"D6", x"A9", x"00", x"85", x"75", x"85",
x"76", x"85", x"77", x"A5", x"B9", x"20", x"22", x"D6",
x"A5", x"AF", x"20", x"22", x"D6", x"A5", x"AE", x"20",
x"22", x"D6", x"A5", x"AD", x"20", x"27", x"D6", x"4C",
x"3C", x"D7", x"D0", x"03", x"4C", x"69", x"D5", x"4A",
x"09", x"80", x"A8", x"90", x"13", x"18", x"A5", x"77",
x"65", x"B6", x"85", x"77", x"A5", x"76", x"65", x"B5",
x"85", x"76", x"A5", x"75", x"65", x"B4", x"85", x"75",
x"66", x"75", x"66", x"76", x"66", x"77", x"66", x"B9",
x"98", x"4A", x"D0", x"DE", x"60", x"85", x"71", x"84",
x"72", x"A0", x"03", x"B1", x"71", x"85", x"B6", x"88",
x"B1", x"71", x"85", x"B5", x"88", x"B1", x"71", x"85",
x"B7", x"45", x"B0", x"85", x"B8", x"A5", x"B7", x"09",
x"80", x"85", x"B4", x"88", x"B1", x"71", x"85", x"B3",
x"A5", x"AC", x"60", x"A5", x"B3", x"F0", x"1F", x"18",
x"65", x"AC", x"90", x"04", x"30", x"1D", x"18", x"2C",
x"10", x"14", x"69", x"80", x"85", x"AC", x"D0", x"03",
x"4C", x"F5", x"D4", x"A5", x"B8", x"85", x"B0", x"60",
x"A5", x"B0", x"49", x"FF", x"30", x"05", x"68", x"68",
x"4C", x"F1", x"D4", x"4C", x"64", x"D5", x"20", x"AB",
x"D7", x"AA", x"F0", x"10", x"18", x"69", x"02", x"B0",
x"F2", x"A2", x"00", x"86", x"B8", x"20", x"7C", x"D4",
x"E6", x"AC", x"F0", x"E7", x"60", x"84", x"20", x"00",
x"00", x"20", x"AB", x"D7", x"A9", x"B5", x"A0", x"D6",
x"A2", x"00", x"86", x"B8", x"20", x"4B", x"D7", x"4C",
x"CD", x"D6", x"20", x"4D", x"D6", x"F0", x"68", x"20",
x"BA", x"D7", x"A9", x"00", x"38", x"E5", x"AC", x"85",
x"AC", x"20", x"73", x"D6", x"E6", x"AC", x"F0", x"BB",
x"A2", x"FD", x"A9", x"01", x"A4", x"B4", x"C4", x"AD",
x"D0", x"0A", x"A4", x"B5", x"C4", x"AE", x"D0", x"04",
x"A4", x"B6", x"C4", x"AF", x"08", x"2A", x"90", x"09",
x"E8", x"95", x"77", x"F0", x"2A", x"10", x"2C", x"A9",
x"01", x"28", x"B0", x"0C", x"06", x"B6", x"26", x"B5",
x"26", x"B4", x"B0", x"E8", x"30", x"D6", x"10", x"E4",
x"A8", x"A5", x"B6", x"E5", x"AF", x"85", x"B6", x"A5",
x"B5", x"E5", x"AE", x"85", x"B5", x"A5", x"B4", x"E5",
x"AD", x"85", x"B4", x"98", x"4C", x"04", x"D7", x"A9",
x"40", x"D0", x"D6", x"0A", x"0A", x"0A", x"0A", x"0A",
x"0A", x"85", x"B9", x"28", x"4C", x"3C", x"D7", x"A2",
x"14", x"4C", x"4E", x"C2", x"A5", x"75", x"85", x"AD",
x"A5", x"76", x"85", x"AE", x"A5", x"77", x"85", x"AF",
x"4C", x"D5", x"D4", x"85", x"71", x"84", x"72", x"A0",
x"03", x"B1", x"71", x"85", x"AF", x"88", x"B1", x"71",
x"85", x"AE", x"88", x"B1", x"71", x"85", x"B0", x"09",
x"80", x"85", x"AD", x"88", x"B1", x"71", x"85", x"AC",
x"84", x"B9", x"60", x"A2", x"A8", x"2C", x"A2", x"A4",
x"A0", x"00", x"F0", x"04", x"A6", x"97", x"A4", x"98",
x"20", x"BA", x"D7", x"86", x"71", x"84", x"72", x"A0",
x"03", x"A5", x"AF", x"91", x"71", x"88", x"A5", x"AE",
x"91", x"71", x"88", x"A5", x"B0", x"09", x"7F", x"25",
x"AD", x"91", x"71", x"88", x"A5", x"AC", x"91", x"71",
x"84", x"B9", x"60", x"A5", x"B7", x"85", x"B0", x"A2",
x"04", x"B5", x"B2", x"95", x"AB", x"CA", x"D0", x"F9",
x"86", x"B9", x"60", x"20", x"BA", x"D7", x"A2", x"05",
x"B5", x"AB", x"95", x"B2", x"CA", x"D0", x"F9", x"86",
x"B9", x"60", x"A5", x"AC", x"F0", x"FB", x"06", x"B9",
x"90", x"F7", x"20", x"59", x"D5", x"D0", x"F2", x"4C",
x"2A", x"D5", x"A5", x"AC", x"F0", x"09", x"A5", x"B0",
x"2A", x"A9", x"FF", x"B0", x"02", x"A9", x"01", x"60",
x"20", x"CA", x"D7", x"85", x"AD", x"A9", x"00", x"85",
x"AE", x"A2", x"88", x"A5", x"AD", x"49", x"FF", x"2A",
x"A9", x"00", x"85", x"AF", x"86", x"AC", x"85", x"B9",
x"85", x"B0", x"4C", x"D0", x"D4", x"46", x"B0", x"60",
x"85", x"73", x"84", x"74", x"A0", x"00", x"B1", x"73",
x"C8", x"AA", x"F0", x"C6", x"B1", x"73", x"45", x"B0",
x"30", x"C4", x"E4", x"AC", x"D0", x"1A", x"B1", x"73",
x"09", x"80", x"C5", x"AD", x"D0", x"12", x"C8", x"B1",
x"73", x"C5", x"AE", x"D0", x"0B", x"C8", x"A9", x"7F",
x"C5", x"B9", x"B1", x"73", x"E5", x"AF", x"F0", x"28",
x"A5", x"B0", x"90", x"02", x"49", x"FF", x"4C", x"D0",
x"D7", x"A5", x"AC", x"F0", x"4A", x"38", x"E9", x"98",
x"24", x"B0", x"10", x"09", x"AA", x"A9", x"FF", x"85",
x"B2", x"20", x"3D", x"D5", x"8A", x"A2", x"AC", x"C9",
x"F9", x"10", x"06", x"20", x"7B", x"D5", x"84", x"B2",
x"60", x"A8", x"A5", x"B0", x"29", x"80", x"46", x"AD",
x"05", x"AD", x"85", x"AD", x"20", x"92", x"D5", x"84",
x"B2", x"60", x"A5", x"AC", x"C9", x"98", x"B0", x"1E",
x"20", x"31", x"D8", x"84", x"B9", x"A5", x"B0", x"84",
x"B0", x"49", x"80", x"2A", x"A9", x"98", x"85", x"AC",
x"A5", x"AF", x"85", x"5B", x"4C", x"D0", x"D4", x"85",
x"AD", x"85", x"AE", x"85", x"AF", x"A8", x"60", x"A0",
x"00", x"A2", x"09", x"94", x"A8", x"CA", x"10", x"FB",
x"90", x"0F", x"C9", x"2D", x"D0", x"04", x"86", x"B1",
x"F0", x"04", x"C9", x"2B", x"D0", x"05", x"20", x"BC",
x"00", x"90", x"5B", x"C9", x"2E", x"F0", x"2E", x"C9",
x"45", x"D0", x"30", x"20", x"BC", x"00", x"90", x"17",
x"C9", x"A4", x"F0", x"0E", x"C9", x"2D", x"F0", x"0A",
x"C9", x"A3", x"F0", x"08", x"C9", x"2B", x"F0", x"04",
x"D0", x"07", x"66", x"AB", x"20", x"BC", x"00", x"90",
x"5C", x"24", x"AB", x"10", x"0E", x"A9", x"00", x"38",
x"E5", x"A9", x"4C", x"DD", x"D8", x"66", x"AA", x"24",
x"AA", x"50", x"C3", x"A5", x"A9", x"38", x"E5", x"A8",
x"85", x"A9", x"F0", x"12", x"10", x"09", x"20", x"B9",
x"D6", x"E6", x"A9", x"D0", x"F9", x"F0", x"07", x"20",
x"9E", x"D6", x"C6", x"A9", x"D0", x"F9", x"A5", x"B1",
x"30", x"01", x"60", x"4C", x"EF", x"DA", x"48", x"24",
x"AA", x"10", x"02", x"E6", x"A8", x"20", x"9E", x"D6",
x"68", x"38", x"E9", x"30", x"20", x"12", x"D9", x"4C",
x"9E", x"D8", x"48", x"20", x"AB", x"D7", x"68", x"20",
x"DB", x"D7", x"A5", x"B7", x"45", x"B0", x"85", x"B8",
x"A6", x"AC", x"4C", x"6F", x"D4", x"A5", x"A9", x"C9",
x"0A", x"90", x"09", x"A9", x"64", x"24", x"AB", x"30",
x"11", x"4C", x"64", x"D5", x"0A", x"0A", x"18", x"65",
x"A9", x"0A", x"18", x"A0", x"00", x"71", x"C3", x"38",
x"E9", x"30", x"85", x"A9", x"4C", x"C4", x"D8", x"91",
x"43", x"4F", x"F8", x"94", x"74", x"23", x"F7", x"94",
x"74", x"24", x"00", x"A9", x"8E", x"A0", x"C1", x"20",
x"6B", x"D9", x"A5", x"88", x"A6", x"87", x"85", x"AD",
x"86", x"AE", x"A2", x"90", x"38", x"20", x"E8", x"D7",
x"20", x"6E", x"D9", x"4C", x"C3", x"C8", x"A0", x"01",
x"A9", x"20", x"24", x"B0", x"10", x"02", x"A9", x"2D",
x"99", x"FF", x"00", x"85", x"B0", x"84", x"BA", x"C8",
x"A9", x"30", x"A6", x"AC", x"D0", x"03", x"4C", x"89",
x"DA", x"A9", x"00", x"E0", x"80", x"F0", x"02", x"B0",
x"09", x"A9", x"4F", x"A0", x"D9", x"20", x"FB", x"D5",
x"A9", x"FA", x"85", x"A8", x"A9", x"4B", x"A0", x"D9",
x"20", x"F8", x"D7", x"F0", x"1E", x"10", x"12", x"A9",
x"47", x"A0", x"D9", x"20", x"F8", x"D7", x"F0", x"02",
x"10", x"0E", x"20", x"9E", x"D6", x"C6", x"A8", x"D0",
x"EE", x"20", x"B9", x"D6", x"E6", x"A8", x"D0", x"DC",
x"20", x"4E", x"D4", x"20", x"31", x"D8", x"A2", x"01",
x"A5", x"A8", x"18", x"69", x"07", x"30", x"09", x"C9",
x"08", x"B0", x"06", x"69", x"FF", x"AA", x"A9", x"02",
x"38", x"E9", x"02", x"85", x"A9", x"86", x"A8", x"8A",
x"F0", x"02", x"10", x"13", x"A4", x"BA", x"A9", x"2E",
x"C8", x"99", x"FF", x"00", x"8A", x"F0", x"06", x"A9",
x"30", x"C8", x"99", x"FF", x"00", x"84", x"BA", x"A0",
x"00", x"A2", x"80", x"A5", x"AF", x"18", x"79", x"9C",
x"DA", x"85", x"AF", x"A5", x"AE", x"79", x"9B", x"DA",
x"85", x"AE", x"A5", x"AD", x"79", x"9A", x"DA", x"85",
x"AD", x"E8", x"B0", x"04", x"10", x"E5", x"30", x"02",
x"30", x"E1", x"8A", x"90", x"04", x"49", x"FF", x"69",
x"0A", x"69", x"2F", x"C8", x"C8", x"C8", x"84", x"95",
x"A4", x"BA", x"C8", x"AA", x"29", x"7F", x"99", x"FF",
x"00", x"C6", x"A8", x"D0", x"06", x"A9", x"2E", x"C8",
x"99", x"FF", x"00", x"84", x"BA", x"A4", x"95", x"8A",
x"49", x"FF", x"29", x"80", x"AA", x"C0", x"12", x"D0",
x"B2", x"A4", x"BA", x"B9", x"FF", x"00", x"88", x"C9",
x"30", x"F0", x"F8", x"C9", x"2E", x"F0", x"01", x"C8",
x"A9", x"2B", x"A6", x"A9", x"F0", x"2E", x"10", x"08",
x"A9", x"00", x"38", x"E5", x"A9", x"AA", x"A9", x"2D",
x"99", x"01", x"01", x"A9", x"45", x"99", x"00", x"01",
x"8A", x"A2", x"2F", x"38", x"E8", x"E9", x"0A", x"B0",
x"FB", x"69", x"3A", x"99", x"03", x"01", x"8A", x"99",
x"02", x"01", x"A9", x"00", x"99", x"04", x"01", x"F0",
x"08", x"99", x"FF", x"00", x"A9", x"00", x"99", x"00",
x"01", x"A9", x"00", x"A0", x"01", x"60", x"80", x"00",
x"00", x"00", x"FE", x"79", x"60", x"00", x"27", x"10",
x"FF", x"FC", x"18", x"00", x"00", x"64", x"FF", x"FF",
x"F6", x"00", x"00", x"01", x"20", x"AB", x"D7", x"A9",
x"96", x"A0", x"DA", x"20", x"4B", x"D7", x"F0", x"63",
x"A5", x"B3", x"D0", x"03", x"4C", x"F3", x"D4", x"A2",
x"9C", x"A0", x"00", x"20", x"78", x"D7", x"A5", x"B7",
x"10", x"0F", x"20", x"62", x"D8", x"A9", x"9C", x"A0",
x"00", x"20", x"F8", x"D7", x"D0", x"03", x"98", x"A4",
x"5B", x"20", x"9D", x"D7", x"98", x"48", x"20", x"BD",
x"D5", x"A9", x"9C", x"A0", x"00", x"20", x"FB", x"D5",
x"20", x"1B", x"DB", x"68", x"4A", x"90", x"0A", x"A5",
x"AC", x"F0", x"06", x"A5", x"B0", x"49", x"FF", x"85",
x"B0", x"60", x"81", x"38", x"AA", x"3B", x"06", x"74",
x"63", x"90", x"8C", x"77", x"23", x"0C", x"AB", x"7A",
x"1E", x"94", x"00", x"7C", x"63", x"42", x"80", x"7E",
x"75", x"FE", x"D0", x"80", x"31", x"72", x"15", x"81",
x"00", x"00", x"00", x"A9", x"FA", x"A0", x"DA", x"20",
x"FB", x"D5", x"A5", x"B9", x"69", x"50", x"90", x"03",
x"20", x"C2", x"D7", x"85", x"A3", x"20", x"AE", x"D7",
x"A5", x"AC", x"C9", x"88", x"90", x"03", x"20", x"90",
x"D6", x"20", x"62", x"D8", x"A5", x"5B", x"18", x"69",
x"81", x"F0", x"F3", x"38", x"E9", x"01", x"48", x"A2",
x"04", x"B5", x"B3", x"B4", x"AC", x"95", x"AC", x"94",
x"B3", x"CA", x"10", x"F5", x"A5", x"A3", x"85", x"B9",
x"20", x"58", x"D4", x"20", x"EF", x"DA", x"A9", x"FE",
x"A0", x"DA", x"20", x"84", x"DB", x"A9", x"00", x"85",
x"B8", x"68", x"20", x"75", x"D6", x"60", x"85", x"BA",
x"84", x"BB", x"20", x"6E", x"D7", x"A9", x"A4", x"20",
x"FB", x"D5", x"20", x"88", x"DB", x"A9", x"A4", x"A0",
x"00", x"4C", x"FB", x"D5", x"85", x"BA", x"84", x"BB",
x"20", x"6B", x"D7", x"B1", x"BA", x"85", x"B1", x"A4",
x"BA", x"C8", x"98", x"D0", x"02", x"E6", x"BB", x"85",
x"BA", x"A4", x"BB", x"20", x"FB", x"D5", x"A5", x"BA",
x"A4", x"BB", x"18", x"69", x"04", x"90", x"01", x"C8",
x"85", x"BA", x"84", x"BB", x"20", x"6C", x"D4", x"A9",
x"A8", x"A0", x"00", x"C6", x"B1", x"D0", x"E4", x"60",
x"98", x"35", x"44", x"7A", x"68", x"28", x"B1", x"46",
x"20", x"CA", x"D7", x"AA", x"30", x"18", x"A9", x"D4",
x"A0", x"00", x"20", x"4B", x"D7", x"8A", x"F0", x"E7",
x"A9", x"B8", x"A0", x"DB", x"20", x"FB", x"D5", x"A9",
x"BC", x"A0", x"DB", x"20", x"6C", x"D4", x"A6", x"AF",
x"A5", x"AD", x"85", x"AF", x"86", x"AD", x"A9", x"00",
x"85", x"B0", x"A5", x"AC", x"85", x"B9", x"A9", x"80",
x"85", x"AC", x"20", x"D5", x"D4", x"A2", x"D4", x"A0",
x"00", x"4C", x"78", x"D7", x"A9", x"78", x"A0", x"DC",
x"20", x"6C", x"D4", x"20", x"AB", x"D7", x"A9", x"7C",
x"A0", x"DC", x"A6", x"B7", x"20", x"C2", x"D6", x"20",
x"AB", x"D7", x"20", x"62", x"D8", x"A9", x"00", x"85",
x"B8", x"20", x"58", x"D4", x"A9", x"80", x"A0", x"DC",
x"20", x"55", x"D4", x"A5", x"B0", x"48", x"10", x"0D",
x"20", x"4E", x"D4", x"A5", x"B0", x"30", x"09", x"A5",
x"63", x"49", x"FF", x"85", x"63", x"20", x"EF", x"DA",
x"A9", x"80", x"A0", x"DC", x"20", x"6C", x"D4", x"68",
x"10", x"03", x"20", x"EF", x"DA", x"A9", x"84", x"A0",
x"DC", x"4C", x"6E", x"DB", x"20", x"6E", x"D7", x"A9",
x"00", x"85", x"63", x"20", x"03", x"DC", x"A2", x"9C",
x"A0", x"00", x"20", x"F9", x"DB", x"A9", x"A4", x"A0",
x"00", x"20", x"4B", x"D7", x"A9", x"00", x"85", x"B0",
x"A5", x"63", x"20", x"74", x"DC", x"A9", x"9C", x"A0",
x"00", x"4C", x"CA", x"D6", x"48", x"4C", x"35", x"DC",
x"81", x"49", x"0F", x"DB", x"83", x"49", x"0F", x"DB",
x"7F", x"00", x"00", x"00", x"04", x"86", x"1E", x"D7",
x"FB", x"87", x"99", x"26", x"65", x"87", x"23", x"34",
x"58", x"86", x"A5", x"5D", x"E1", x"83", x"49", x"0F",
x"DB", x"A5", x"B0", x"48", x"10", x"03", x"20", x"EF",
x"DA", x"A5", x"AC", x"48", x"C9", x"81", x"90", x"07",
x"A9", x"9C", x"A0", x"D5", x"20", x"CA", x"D6", x"A9",
x"C9", x"A0", x"DC", x"20", x"6E", x"DB", x"68", x"C9",
x"81", x"90", x"07", x"A9", x"78", x"A0", x"DC", x"20",
x"55", x"D4", x"68", x"10", x"03", x"4C", x"EF", x"DA",
x"60", x"08", x"78", x"3A", x"C5", x"37", x"7B", x"83",
x"A2", x"5C", x"7C", x"2E", x"DD", x"4D", x"7D", x"99",
x"B0", x"1E", x"7D", x"59", x"ED", x"24", x"7E", x"91",
x"72", x"00", x"7E", x"4C", x"B9", x"73", x"7F", x"AA",
x"AA", x"53", x"81", x"00", x"00", x"00", x"E6", x"C3",
x"D0", x"02", x"E6", x"C4", x"AD", x"DD", x"DD", x"C9",
x"3A", x"B0", x"0A", x"C9", x"20", x"F0", x"EF", x"38",
x"E9", x"30", x"38", x"E9", x"D0", x"60", x"80", x"4F",
x"C7", x"52", x"A9", x"39", x"A0", x"DE", x"20", x"C3",
x"C8", x"A2", x"FF", x"86", x"88", x"9A", x"A9", x"11",
x"A0", x"DD", x"85", x"01", x"84", x"02", x"85", x"04",
x"84", x"05", x"A9", x"05", x"A0", x"CE", x"85", x"06",
x"84", x"07", x"A9", x"C1", x"A0", x"CF", x"85", x"08",
x"84", x"09", x"A9", x"4C", x"85", x"00", x"85", x"03",
x"85", x"A1", x"85", x"0A", x"A9", x"88", x"A0", x"CE",
x"85", x"0B", x"84", x"0C", x"A9", x"3F", x"85", x"0F",
x"A9", x"38", x"85", x"10", x"A2", x"1C", x"BD", x"ED",
x"DC", x"95", x"BB", x"CA", x"D0", x"F8", x"8A", x"85",
x"B2", x"85", x"67", x"85", x"0D", x"85", x"0E", x"48",
x"85", x"64", x"A9", x"03", x"85", x"A0", x"A9", x"2C",
x"85", x"12", x"20", x"6C", x"C8", x"A2", x"68", x"86",
x"65", x"A9", x"5A", x"A0", x"DE", x"20", x"C3", x"C8",
x"20", x"46", x"C9", x"86", x"C3", x"84", x"C4", x"20",
x"BC", x"00", x"C9", x"41", x"F0", x"84", x"A8", x"D0",
x"21", x"A9", x"00", x"A0", x"04", x"85", x"11", x"84",
x"12", x"A0", x"00", x"E6", x"11", x"D0", x"02", x"E6",
x"12", x"4C", x"A3", x"DE", x"EA", x"D1", x"11", x"D0",
x"15", x"0A", x"91", x"11", x"D1", x"11", x"F0", x"EB",
x"D0", x"0C", x"20", x"C2", x"00", x"20", x"7F", x"C7",
x"A8", x"F0", x"03", x"4C", x"0C", x"CC", x"A5", x"11",
x"A4", x"12", x"85", x"85", x"84", x"86", x"85", x"81",
x"84", x"82", x"A9", x"66", x"A0", x"DE", x"20", x"C3",
x"C8", x"20", x"46", x"C9", x"86", x"C3", x"84", x"C4",
x"20", x"BC", x"00", x"A8", x"F0", x"1C", x"20", x"7F",
x"C7", x"A5", x"12", x"D0", x"E5", x"A5", x"11", x"C9",
x"10", x"90", x"DF", x"85", x"0F", x"E9", x"0E", x"B0",
x"FC", x"49", x"FF", x"E9", x"0C", x"18", x"65", x"0F",
x"85", x"10", x"A2", x"00", x"A0", x"04", x"86", x"79",
x"84", x"7A", x"A0", x"00", x"98", x"91", x"79", x"E6",
x"79", x"D0", x"02", x"E6", x"7A", x"A5", x"79", x"A4",
x"7A", x"20", x"1F", x"C2", x"20", x"6C", x"C8", x"A5",
x"85", x"38", x"E5", x"79", x"AA", x"A5", x"86", x"E5",
x"7A", x"20", x"5E", x"D9", x"A9", x"75", x"A0", x"DE",
x"20", x"C3", x"C8", x"A9", x"C3", x"A0", x"C8", x"85",
x"04", x"84", x"05", x"20", x"63", x"C4", x"A9", x"74",
x"A0", x"C2", x"85", x"01", x"84", x"02", x"6C", x"01",
x"00", x"42", x"41", x"53", x"49", x"43", x"2D", x"50",
x"52", x"49", x"56", x"52", x"45", x"4D", x"45", x"4E",
x"41", x"20", x"56", x"45", x"52", x"5A", x"49", x"4A",
x"41", x"20", x"38", x"34", x"30", x"31", x"32", x"34",
x"0C", x"00", x"20", x"4D", x"45", x"4D", x"4F", x"52",
x"49", x"4A", x"41", x"20", x"20", x"00", x"44", x"55",
x"4C", x"4A", x"49", x"4E", x"41", x"20", x"4C", x"49",
x"4E", x"49", x"4A", x"45", x"00", x"20", x"4C", x"4F",
x"4B", x"41", x"43", x"49", x"4A", x"41", x"0D", x"0A",
x"00", x"20", x"FC", x"D3", x"A5", x"11", x"85", x"E4",
x"86", x"E5", x"4C", x"8B", x"FE", x"20", x"FC", x"D3",
x"A5", x"11", x"85", x"E2", x"86", x"E3", x"4C", x"69",
x"FE", x"20", x"FC", x"D3", x"A5", x"11", x"85", x"E2",
x"86", x"E3", x"60", x"A5", x"12", x"C9", x"60", x"F0",
x"07", x"A9", x"92", x"91", x"11", x"4C", x"9D", x"DD",
x"4C", x"B6", x"DD", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			data <= romData(conv_integer(addr));
		end if;
	end process;
end architecture;

