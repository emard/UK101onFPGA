library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity rom_crt is
	port (
		clk: in std_logic;
		addr: in std_logic_vector(12 downto 0);
		data: out std_logic_vector(7 downto 0)
	);
end entity;

architecture Behavioral of rom_crt is
	type romDef is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant romData: romDef := (
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"08", x"08", x"08", x"08", x"08", x"00", x"08", x"00",
x"14", x"14", x"00", x"00", x"00", x"00", x"00", x"00",
x"28", x"28", x"7C", x"28", x"7C", x"28", x"28", x"00",
x"10", x"78", x"14", x"38", x"50", x"3C", x"10", x"00",
x"46", x"26", x"10", x"08", x"64", x"62", x"00", x"00",
x"08", x"14", x"14", x"0C", x"52", x"22", x"5C", x"00",
x"20", x"10", x"08", x"00", x"00", x"00", x"00", x"00",
x"20", x"10", x"08", x"08", x"08", x"10", x"20", x"00",
x"04", x"08", x"10", x"10", x"10", x"08", x"04", x"00",
x"00", x"10", x"54", x"38", x"54", x"10", x"00", x"00",
x"00", x"10", x"10", x"7C", x"10", x"10", x"00", x"00",
x"00", x"00", x"00", x"00", x"18", x"18", x"04", x"00",
x"00", x"00", x"00", x"7C", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00",
x"00", x"40", x"20", x"10", x"08", x"04", x"00", x"00",
x"38", x"44", x"64", x"54", x"4C", x"44", x"38", x"00",
x"10", x"18", x"10", x"10", x"10", x"10", x"38", x"00",
x"38", x"44", x"40", x"20", x"18", x"04", x"7C", x"00",
x"7C", x"20", x"10", x"20", x"40", x"44", x"38", x"00",
x"20", x"30", x"28", x"24", x"7C", x"20", x"20", x"00",
x"7C", x"04", x"3C", x"40", x"40", x"44", x"38", x"00",
x"30", x"08", x"04", x"3C", x"44", x"44", x"38", x"00",
x"7C", x"40", x"20", x"10", x"08", x"08", x"08", x"00",
x"38", x"44", x"44", x"38", x"44", x"44", x"38", x"00",
x"38", x"44", x"44", x"78", x"40", x"20", x"18", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"04", x"00",
x"20", x"10", x"08", x"04", x"08", x"10", x"20", x"00",
x"00", x"00", x"7C", x"00", x"7C", x"00", x"00", x"00",
x"04", x"08", x"10", x"20", x"10", x"08", x"04", x"00",
x"1C", x"22", x"20", x"18", x"08", x"00", x"08", x"00",
x"38", x"44", x"74", x"54", x"74", x"04", x"78", x"00",
x"38", x"44", x"44", x"7C", x"44", x"44", x"44", x"00",
x"3C", x"48", x"48", x"38", x"48", x"48", x"3C", x"00",
x"38", x"44", x"04", x"04", x"04", x"44", x"38", x"00",
x"3C", x"48", x"48", x"48", x"48", x"48", x"3C", x"00",
x"7C", x"04", x"04", x"1C", x"04", x"04", x"7C", x"00",
x"7C", x"04", x"04", x"1C", x"04", x"04", x"04", x"00",
x"38", x"44", x"04", x"04", x"74", x"44", x"78", x"00",
x"44", x"44", x"44", x"7C", x"44", x"44", x"44", x"00",
x"38", x"10", x"10", x"10", x"10", x"10", x"38", x"00",
x"70", x"20", x"20", x"20", x"20", x"24", x"18", x"00",
x"44", x"24", x"14", x"0C", x"14", x"24", x"44", x"00",
x"04", x"04", x"04", x"04", x"04", x"04", x"7C", x"00",
x"44", x"6C", x"54", x"54", x"44", x"44", x"44", x"00",
x"44", x"44", x"4C", x"54", x"64", x"44", x"44", x"00",
x"38", x"44", x"44", x"44", x"44", x"44", x"38", x"00",
x"3C", x"44", x"44", x"3C", x"04", x"04", x"04", x"00",
x"38", x"44", x"44", x"44", x"54", x"24", x"58", x"00",
x"3C", x"44", x"44", x"3C", x"14", x"24", x"44", x"00",
x"38", x"44", x"08", x"10", x"20", x"44", x"38", x"00",
x"7C", x"10", x"10", x"10", x"10", x"10", x"10", x"00",
x"44", x"44", x"44", x"44", x"44", x"44", x"38", x"00",
x"44", x"44", x"44", x"44", x"44", x"28", x"10", x"00",
x"44", x"44", x"44", x"54", x"54", x"54", x"28", x"00",
x"44", x"44", x"28", x"10", x"28", x"44", x"44", x"00",
x"44", x"44", x"44", x"28", x"10", x"10", x"10", x"00",
x"7C", x"40", x"20", x"10", x"08", x"04", x"7C", x"00",
x"28", x"38", x"44", x"04", x"04", x"44", x"38", x"00",
x"20", x"38", x"44", x"04", x"04", x"44", x"38", x"00",
x"3C", x"48", x"48", x"5C", x"48", x"48", x"3C", x"00",
x"28", x"38", x"44", x"08", x"30", x"44", x"38", x"00",
x"28", x"7C", x"40", x"20", x"10", x"08", x"7C", x"00",
x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00",
x"00", x"18", x"20", x"38", x"24", x"38", x"00", x"00",
x"04", x"04", x"1C", x"24", x"24", x"1C", x"00", x"00",
x"00", x"38", x"04", x"04", x"04", x"38", x"00", x"00",
x"20", x"20", x"38", x"24", x"24", x"38", x"00", x"00",
x"00", x"18", x"24", x"1C", x"04", x"18", x"00", x"00",
x"10", x"28", x"08", x"1C", x"08", x"08", x"08", x"00",
x"00", x"38", x"24", x"24", x"38", x"20", x"18", x"00",
x"04", x"04", x"1C", x"24", x"24", x"24", x"00", x"00",
x"10", x"00", x"18", x"10", x"10", x"38", x"00", x"00",
x"10", x"00", x"18", x"10", x"10", x"14", x"08", x"00",
x"04", x"04", x"14", x"0C", x"14", x"24", x"00", x"00",
x"18", x"10", x"10", x"10", x"10", x"38", x"00", x"00",
x"00", x"2C", x"54", x"54", x"54", x"54", x"00", x"00",
x"00", x"1C", x"24", x"24", x"24", x"24", x"00", x"00",
x"00", x"18", x"24", x"24", x"24", x"18", x"00", x"00",
x"00", x"1C", x"24", x"24", x"1C", x"04", x"04", x"00",
x"00", x"1C", x"12", x"12", x"1C", x"10", x"78", x"00",
x"00", x"34", x"0C", x"04", x"04", x"04", x"00", x"00",
x"00", x"38", x"04", x"18", x"20", x"1C", x"00", x"00",
x"10", x"38", x"10", x"10", x"10", x"20", x"00", x"00",
x"00", x"24", x"24", x"24", x"24", x"38", x"00", x"00",
x"00", x"44", x"44", x"44", x"28", x"10", x"00", x"00",
x"00", x"44", x"44", x"54", x"54", x"28", x"00", x"00",
x"00", x"44", x"28", x"10", x"28", x"44", x"00", x"00",
x"00", x"24", x"24", x"24", x"38", x"20", x"18", x"00",
x"00", x"3C", x"20", x"10", x"08", x"3C", x"00", x"00",
x"38", x"00", x"38", x"04", x"04", x"38", x"00", x"00",
x"20", x"00", x"38", x"04", x"04", x"38", x"00", x"00",
x"20", x"70", x"20", x"38", x"24", x"38", x"00", x"00",
x"28", x"38", x"04", x"18", x"20", x"1C", x"00", x"00",
x"38", x"00", x"3C", x"10", x"08", x"3C", x"00", x"00",
x"09", x"0A", x"0B", x"08", x"14", x"13", x"12", x"11",
x"36", x"74", x"7A", x"72", x"37", x"75", x"69", x"6F",
x"31", x"77", x"71", x"65", x"6D", x"6B", x"6A", x"6C",
x"79", x"73", x"61", x"64", x"6E", x"67", x"68", x"66",
x"3A", x"7F", x"7C", x"7B", x"3B", x"7E", x"7D", x"70",
x"00", x"0D", x"00", x"20", x"34", x"35", x"39", x"38",
x"33", x"32", x"2E", x"2C", x"63", x"78", x"76", x"62",
x"60", x"2F", x"30", x"2D", x"87", x"FC", x"87", x"FA",
x"87", x"F6", x"87", x"EE", x"87", x"DE", x"87", x"BE",
x"87", x"7E", x"86", x"FE", x"85", x"FE", x"83", x"FE",
x"85", x"FC", x"8A", x"48", x"98", x"48", x"A5", x"FC",
x"A8", x"2A", x"2A", x"2A", x"2A", x"29", x"03", x"AA",
x"BD", x"00", x"02", x"D0", x"05", x"BD", x"04", x"02",
x"F0", x"24", x"85", x"F1", x"98", x"0A", x"0A", x"0A",
x"85", x"F0", x"A0", x"07", x"B1", x"F0", x"84", x"FA",
x"A4", x"E9", x"24", x"FC", x"10", x"02", x"49", x"FF",
x"91", x"E6", x"A5", x"E6", x"38", x"E9", x"20", x"85",
x"E6", x"A4", x"FA", x"88", x"10", x"E6", x"68", x"A8",
x"68", x"AA", x"A5", x"FC", x"60", x"A6", x"EA", x"86",
x"E8", x"A4", x"EC", x"84", x"E9", x"A9", x"E0", x"85",
x"E6", x"A5", x"E8", x"20", x"9E", x"EE", x"60", x"EA",
x"EA", x"EA", x"A6", x"EB", x"18", x"90", x"05", x"20",
x"95", x"E3", x"A4", x"EC", x"20", x"AD", x"E4", x"C4",
x"ED", x"C8", x"90", x"F8", x"E4", x"EB", x"B0", x"15",
x"E8", x"E6", x"E7", x"90", x"ED", x"C6", x"E9", x"C4",
x"EC", x"D0", x"0D", x"A4", x"ED", x"84", x"E9", x"E4",
x"EA", x"F0", x"05", x"C6", x"E8", x"20", x"9D", x"E3",
x"68", x"A8", x"68", x"AA", x"A5", x"FC", x"60", x"85",
x"FC", x"8A", x"48", x"98", x"48", x"A5", x"FC", x"A6",
x"E8", x"A4", x"E9", x"C9", x"20", x"B0", x"39", x"2C",
x"08", x"02", x"30", x"34", x"4C", x"B0", x"EE", x"EA",
x"C9", x"0C", x"F0", x"B3", x"C9", x"06", x"F0", x"B4",
x"C9", x"08", x"F0", x"C1", x"C9", x"0B", x"F0", x"C7",
x"C9", x"09", x"F0", x"1F", x"C9", x"0A", x"F0", x"25",
x"C9", x"0D", x"F0", x"6A", x"C9", x"04", x"D0", x"06",
x"20", x"95", x"E3", x"4C", x"D8", x"E3", x"C9", x"07",
x"D0", x"B6", x"20", x"F4", x"E4", x"4C", x"D8", x"E3",
x"20", x"50", x"E3", x"E6", x"E9", x"C4", x"ED", x"90",
x"A7", x"A4", x"EC", x"84", x"E9", x"E6", x"E8", x"E4",
x"EB", x"90", x"9A", x"C6", x"E8", x"A5", x"EA", x"20",
x"A3", x"E3", x"A5", x"E6", x"18", x"90", x"13", x"E6",
x"E7", x"A4", x"EC", x"B1", x"E6", x"91", x"EE", x"C4",
x"ED", x"C8", x"90", x"F7", x"A5", x"E6", x"E9", x"20",
x"85", x"E6", x"85", x"EE", x"B0", x"EB", x"A5", x"E7",
x"85", x"EF", x"38", x"E9", x"60", x"C5", x"EB", x"90",
x"DE", x"4C", x"B2", x"E3", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"20", x"0F",
x"E6", x"F0", x"1C", x"A0", x"09", x"88", x"F0", x"17",
x"A2", x"FF", x"20", x"E3", x"E4", x"20", x"0F", x"E6",
x"D0", x"F3", x"A4", x"E9", x"20", x"C2", x"E4", x"20",
x"0F", x"E6", x"F0", x"FB", x"20", x"C2", x"E4", x"A6",
x"E8", x"AD", x"09", x"02", x"D0", x"8B", x"A4", x"EC",
x"84", x"E9", x"4C", x"D8", x"E3", x"86", x"FB", x"A2",
x"08", x"A9", x"00", x"91", x"E6", x"A5", x"E6", x"38",
x"E9", x"20", x"85", x"E6", x"CA", x"D0", x"F2", x"A6",
x"FB", x"60", x"86", x"FB", x"A2", x"08", x"B1", x"E6",
x"49", x"FF", x"91", x"E6", x"A5", x"E6", x"38", x"E9",
x"20", x"85", x"E6", x"CA", x"D0", x"F0", x"A6", x"FB",
x"60", x"48", x"98", x"A0", x"BB", x"88", x"D0", x"FD",
x"A8", x"68", x"60", x"20", x"D9", x"E4", x"CA", x"D0",
x"FA", x"60", x"8E", x"00", x"88", x"20", x"D9", x"E4",
x"CA", x"D0", x"F7", x"60", x"48", x"8A", x"A2", x"70",
x"20", x"EA", x"E4", x"AA", x"68", x"60", x"FF", x"FF",
x"8A", x"48", x"98", x"48", x"A4", x"E9", x"B1", x"E6",
x"48", x"A4", x"E9", x"B1", x"E6", x"49", x"FF", x"91",
x"E6", x"A0", x"00", x"88", x"F0", x"F3", x"20", x"B0",
x"E5", x"90", x"F8", x"85", x"FC", x"F0", x"F4", x"A2",
x"0A", x"20", x"E3", x"E4", x"20", x"B0", x"E5", x"90",
x"EA", x"C5", x"FC", x"D0", x"E6", x"A4", x"E9", x"68",
x"91", x"E6", x"AD", x"0B", x"02", x"F0", x"05", x"A2",
x"0F", x"20", x"EA", x"E4", x"A2", x"04", x"20", x"E3",
x"E4", x"20", x"B0", x"E5", x"90", x"12", x"C5", x"FC",
x"D0", x"0E", x"AE", x"0C", x"02", x"F0", x"ED", x"CE",
x"0C", x"02", x"D0", x"E8", x"A2", x"20", x"D0", x"07",
x"AE", x"0C", x"02", x"F0", x"05", x"A2", x"FF", x"8E",
x"0C", x"02", x"AD", x"FB", x"87", x"29", x"20", x"0A",
x"85", x"FA", x"AD", x"FD", x"87", x"29", x"20", x"05",
x"FA", x"0A", x"85", x"FA", x"A5", x"FC", x"C9", x"21",
x"90", x"2D", x"C9", x"60", x"B0", x"0F", x"2C", x"0E",
x"02", x"10", x"02", x"09", x"80", x"A4", x"FA", x"30",
x"1E", x"49", x"10", x"D0", x"1A", x"F0", x"05", x"2C",
x"0D", x"02", x"10", x"04", x"A4", x"FA", x"30", x"02",
x"49", x"20", x"2C", x"0E", x"02", x"10", x"02", x"09",
x"80", x"24", x"FA", x"70", x"02", x"29", x"1F", x"85",
x"FC", x"68", x"A8", x"68", x"AA", x"A5", x"FC", x"60",
x"8A", x"48", x"98", x"48", x"A2", x"14", x"CA", x"CA",
x"30", x"2D", x"BD", x"3C", x"E3", x"85", x"F1", x"BD",
x"3D", x"E3", x"85", x"F0", x"20", x"F9", x"E5", x"90",
x"ED", x"C0", x"00", x"D0", x"21", x"0A", x"B0", x"09",
x"C8", x"0A", x"B0", x"05", x"C8", x"0A", x"B0", x"01",
x"C8", x"8A", x"0A", x"84", x"FA", x"18", x"65", x"FA",
x"AA", x"BD", x"00", x"E3", x"85", x"FA", x"38", x"68",
x"A8", x"68", x"AA", x"A5", x"FA", x"60", x"29", x"10",
x"D0", x"01", x"88", x"8A", x"18", x"69", x"28", x"D0",
x"E2", x"38", x"A0", x"00", x"B1", x"F0", x"09", x"0F",
x"49", x"FF", x"D0", x"0A", x"C8", x"B1", x"F0", x"09",
x"CF", x"49", x"FF", x"D0", x"01", x"18", x"60", x"AD",
x"00", x"80", x"09", x"0F", x"49", x"FF", x"D0", x"07",
x"AD", x"01", x"80", x"09", x"CF", x"49", x"FF", x"60",
x"20", x"33", x"E6", x"C9", x"57", x"D0", x"03", x"4C",
x"74", x"C2", x"C9", x"43", x"D0", x"03", x"4C", x"11",
x"DD", x"60", x"E8", x"BD", x"80", x"02", x"C9", x"20",
x"F0", x"F8", x"60", x"85", x"F3", x"84", x"F2", x"98",
x"48", x"A0", x"00", x"B1", x"F2", x"C9", x"04", x"F0",
x"0B", x"20", x"F1", x"FF", x"E6", x"F2", x"D0", x"F3",
x"E6", x"F3", x"D0", x"EF", x"68", x"A8", x"60", x"A2",
x"00", x"8A", x"F0", x"01", x"CA", x"20", x"EE", x"FF",
x"9D", x"80", x"02", x"C9", x"0D", x"F0", x"1B", x"C9",
x"08", x"F0", x"EE", x"C9", x"18", x"F0", x"0D", x"C9",
x"20", x"90", x"EA", x"E8", x"10", x"E7", x"20", x"F4",
x"E4", x"38", x"B0", x"E0", x"A9", x"0D", x"A2", x"00",
x"F0", x"DE", x"60", x"FF", x"0D", x"0A", x"00", x"00",
x"00", x"00", x"2A", x"04", x"E0", x"2F", x"00", x"00",
x"00", x"00", x"E0", x"60", x"00", x"00", x"00", x"1F",
x"00", x"1F", x"E0", x"20", x"00", x"00", x"00", x"00",
x"00", x"E0", x"E1", x"E2", x"00", x"00", x"00", x"00",
x"FF", x"00", x"00", x"00", x"00", x"FF", x"FD", x"2A",
x"FF", x"FF", x"1C", x"E7", x"62", x"E7", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"20", x"E6", x"FD", x"E8", x"06", x"E9", x"0E", x"E9",
x"D0", x"EA", x"09", x"EB", x"48", x"EB", x"6A", x"EB",
x"AB", x"EB", x"80", x"EC", x"F6", x"EE", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"42", x"4A", x"55", x"45", x"43", x"51", x"46", x"4D",
x"41", x"58", x"50", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"20", x"00", x"E5", x"C9",
x"11", x"90", x"09", x"C9", x"14", x"B0", x"05", x"20",
x"34", x"E7", x"A9", x"00", x"2C", x"0F", x"02", x"30",
x"30", x"4C", x"F1", x"FF", x"C9", x"12", x"90", x"21",
x"F0", x"16", x"C9", x"13", x"B0", x"09", x"AD", x"0B",
x"02", x"49", x"FF", x"8D", x"0B", x"02", x"60", x"AD",
x"0E", x"02", x"49", x"FF", x"8D", x"0E", x"02", x"60",
x"AD", x"10", x"02", x"49", x"FF", x"8D", x"10", x"02",
x"60", x"AD", x"0D", x"02", x"49", x"FF", x"8D", x"0D",
x"02", x"60", x"20", x"DF", x"E3", x"2C", x"10", x"02",
x"10", x"F7", x"4C", x"E9", x"EE", x"EA", x"EA", x"BA",
x"BD", x"03", x"01", x"A2", x"09", x"18", x"2A", x"6A",
x"B0", x"05", x"8D", x"00", x"98", x"90", x"07", x"29",
x"FF", x"30", x"03", x"8D", x"00", x"90", x"AC", x"13",
x"02", x"20", x"B8", x"E7", x"CA", x"30", x"06", x"D0",
x"E6", x"09", x"01", x"D0", x"E2", x"68", x"A8", x"68",
x"AA", x"68", x"60", x"FF", x"FF", x"FF", x"FF", x"A0",
x"00", x"8C", x"00", x"98", x"8C", x"00", x"90", x"2C",
x"FF", x"87", x"10", x"03", x"C8", x"D0", x"F8", x"88",
x"84", x"F4", x"60", x"AE", x"2A", x"0A", x"04", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"88", x"D0",
x"F6", x"60", x"FF", x"48", x"10", x"05", x"38", x"90",
x"02", x"49", x"80", x"0A", x"D0", x"F9", x"68", x"60",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"48", x"A9", x"20", x"20",
x"F1", x"FF", x"68", x"60", x"A2", x"03", x"20", x"DC",
x"E7", x"CA", x"D0", x"FA", x"60", x"C9", x"0A", x"90",
x"02", x"69", x"06", x"69", x"30", x"60", x"A9", x"0D",
x"20", x"F1", x"FF", x"A9", x"0A", x"4C", x"F1", x"FF",
x"20", x"DC", x"E7", x"48", x"4A", x"4A", x"4A", x"4A",
x"20", x"ED", x"E7", x"20", x"F1", x"FF", x"68", x"29",
x"0F", x"20", x"ED", x"E7", x"4C", x"F1", x"FF", x"20",
x"DC", x"E7", x"A5", x"FF", x"20", x"03", x"E8", x"A5",
x"FE", x"4C", x"03", x"E8", x"20", x"33", x"E6", x"BD",
x"80", x"02", x"E8", x"C9", x"30", x"90", x"0F", x"E9",
x"30", x"C9", x"0A", x"90", x"0A", x"C9", x"11", x"90",
x"05", x"E9", x"07", x"C9", x"10", x"60", x"38", x"60",
x"20", x"27", x"E8", x"90", x"06", x"60", x"20", x"24",
x"E8", x"B0", x"0F", x"0A", x"0A", x"0A", x"0A", x"85",
x"FC", x"20", x"27", x"E8", x"B0", x"04", x"05", x"FC",
x"85", x"FC", x"60", x"20", x"46", x"E8", x"B0", x"07",
x"85", x"F7", x"20", x"40", x"E8", x"85", x"F6", x"60",
x"20", x"7D", x"E8", x"B0", x"1D", x"20", x"92", x"E8",
x"B0", x"18", x"4C", x"5B", x"E8", x"20", x"7D", x"E8",
x"B0", x"10", x"4C", x"5B", x"E8", x"20", x"5B", x"E8",
x"B0", x"08", x"A5", x"F6", x"85", x"FE", x"A5", x"F7",
x"85", x"FF", x"60", x"E6", x"FE", x"D0", x"02", x"E6",
x"FF", x"60", x"20", x"5B", x"E8", x"B0", x"08", x"A5",
x"F6", x"85", x"F4", x"A5", x"F7", x"85", x"F5", x"60",
x"E6", x"F4", x"D0", x"02", x"E6", x"F5", x"60", x"18",
x"A5", x"FE", x"65", x"F6", x"85", x"FE", x"A5", x"FF",
x"65", x"F7", x"85", x"FF", x"60", x"38", x"A5", x"FE",
x"E5", x"F4", x"85", x"FE", x"A5", x"FF", x"E5", x"F5",
x"85", x"FF", x"60", x"38", x"A5", x"F6", x"E5", x"F4",
x"A5", x"F7", x"E5", x"F5", x"60", x"38", x"A5", x"FE",
x"E5", x"F4", x"A5", x"FF", x"E5", x"F5", x"60", x"18",
x"A5", x"F6", x"E9", x"00", x"85", x"F6", x"A5", x"F7",
x"E9", x"00", x"85", x"F7", x"60", x"18", x"A5", x"FE",
x"E9", x"00", x"85", x"FE", x"A5", x"FF", x"E9", x"00",
x"85", x"FF", x"60", x"38", x"A5", x"FE", x"E5", x"F6",
x"A5", x"FF", x"E5", x"F7", x"60", x"20", x"5B", x"E8",
x"B0", x"2C", x"68", x"68", x"90", x"05", x"20", x"5B",
x"E8", x"B0", x"23", x"6C", x"F6", x"00", x"20", x"75",
x"E8", x"B0", x"1B", x"A0", x"00", x"20", x"F6", x"E7",
x"20", x"17", x"E8", x"A2", x"09", x"CA", x"F0", x"F5",
x"B1", x"FE", x"20", x"00", x"E8", x"20", x"F3", x"E8",
x"20", x"8B", x"E8", x"90", x"F0", x"18", x"60", x"FF",
x"00", x"90", x"6D", x"65", x"69", x"7D", x"79", x"61",
x"71", x"75", x"D0", x"2D", x"25", x"29", x"3D", x"39",
x"21", x"31", x"35", x"30", x"0A", x"0E", x"06", x"1E",
x"16", x"08", x"90", x"08", x"B0", x"88", x"F0", x"48",
x"2C", x"24", x"C8", x"30", x"C8", x"D0", x"28", x"10",
x"28", x"00", x"A8", x"50", x"A8", x"70", x"D8", x"18",
x"D8", x"D8", x"D8", x"58", x"D8", x"B8", x"D8", x"CD",
x"C5", x"C9", x"DD", x"D9", x"C1", x"D1", x"D5", x"38",
x"EC", x"E4", x"E0", x"38", x"CC", x"C4", x"C0", x"84",
x"CE", x"C6", x"DE", x"D6", x"84", x"CA", x"84", x"88",
x"D4", x"4D", x"45", x"49", x"5D", x"59", x"41", x"51",
x"55", x"D2", x"EE", x"E6", x"FE", x"F6", x"D2", x"E8",
x"D2", x"C8", x"CA", x"4C", x"6C", x"2A", x"20", x"86",
x"AD", x"A5", x"A9", x"BD", x"B9", x"A1", x"B1", x"B5",
x"86", x"AE", x"A6", x"A2", x"BE", x"B6", x"86", x"AC",
x"A4", x"A0", x"BC", x"B4", x"26", x"4A", x"4E", x"46",
x"5E", x"56", x"CE", x"EA", x"3E", x"0D", x"05", x"09",
x"1D", x"19", x"01", x"11", x"15", x"41", x"48", x"41",
x"08", x"C1", x"68", x"C1", x"28", x"C9", x"2A", x"2E",
x"26", x"3E", x"36", x"C9", x"6A", x"6E", x"66", x"7E",
x"76", x"A9", x"40", x"A9", x"60", x"19", x"ED", x"E5",
x"E9", x"FD", x"F9", x"E1", x"F1", x"F5", x"99", x"38",
x"99", x"F8", x"99", x"78", x"B9", x"8D", x"85", x"9D",
x"99", x"81", x"91", x"95", x"B9", x"8E", x"86", x"96",
x"B9", x"8C", x"84", x"94", x"05", x"AA", x"05", x"A8",
x"25", x"BA", x"65", x"8A", x"65", x"9A", x"65", x"98",
x"00", x"60", x"82", x"81", x"C1", x"8A", x"86", x"99",
x"95", x"89", x"11", x"82", x"81", x"C1", x"8A", x"86",
x"99", x"95", x"89", x"1B", x"80", x"82", x"81", x"8A",
x"89", x"63", x"A1", x"67", x"A1", x"46", x"A1", x"16",
x"82", x"81", x"4A", x"A1", x"51", x"A1", x"18", x"A1",
x"69", x"80", x"61", x"A1", x"65", x"A1", x"60", x"80",
x"10", x"80", x"48", x"80", x"34", x"80", x"06", x"82",
x"81", x"C1", x"8A", x"86", x"99", x"95", x"89", x"0C",
x"82", x"81", x"C1", x"4C", x"82", x"81", x"C1", x"62",
x"82", x"81", x"8A", x"89", x"0E", x"80", x"4E", x"80",
x"27", x"82", x"81", x"C1", x"8A", x"86", x"99", x"95",
x"89", x"61", x"82", x"81", x"8A", x"89", x"0D", x"80",
x"4D", x"80", x"06", x"82", x"92", x"27", x"82", x"40",
x"82", x"81", x"C1", x"8A", x"86", x"99", x"95", x"89",
x"0C", x"82", x"81", x"C1", x"86", x"85", x"4C", x"82",
x"81", x"C1", x"8A", x"89", x"27", x"80", x"82", x"81",
x"8A", x"89", x"07", x"80", x"41", x"82", x"81", x"C1",
x"8A", x"86", x"99", x"95", x"89", x"40", x"80", x"04",
x"80", x"40", x"80", x"04", x"80", x"1B", x"80", x"82",
x"81", x"8A", x"89", x"27", x"80", x"82", x"81", x"8A",
x"89", x"48", x"80", x"64", x"80", x"61", x"82", x"81",
x"C1", x"8A", x"86", x"99", x"95", x"89", x"62", x"80",
x"12", x"80", x"4A", x"80", x"40", x"82", x"81", x"8A",
x"86", x"99", x"95", x"89", x"0C", x"82", x"81", x"85",
x"4C", x"82", x"81", x"89", x"0E", x"80", x"4E", x"80",
x"0F", x"80", x"40", x"80", x"64", x"80", x"42", x"80",
x"20", x"75", x"E8", x"B0", x"33", x"A2", x"00", x"86",
x"F4", x"86", x"F5", x"A0", x"00", x"8A", x"71", x"FE",
x"AA", x"90", x"06", x"E6", x"F4", x"D0", x"02", x"E6",
x"F5", x"20", x"F3", x"E8", x"20", x"8B", x"E8", x"90",
x"EC", x"20", x"F6", x"E7", x"A9", x"3D", x"20", x"F1",
x"FF", x"A5", x"F5", x"20", x"00", x"E8", x"A5", x"F4",
x"20", x"00", x"E8", x"8A", x"20", x"00", x"E8", x"18",
x"60", x"20", x"68", x"E8", x"B0", x"25", x"20", x"C3",
x"E8", x"90", x"33", x"A0", x"00", x"20", x"CD", x"E8",
x"90", x"1A", x"20", x"B5", x"E8", x"20", x"A7", x"E8",
x"B0", x"11", x"B1", x"F6", x"91", x"FE", x"20", x"D7",
x"E8", x"90", x"08", x"20", x"E5", x"E8", x"20", x"C3",
x"E8", x"B0", x"EF", x"60", x"B1", x"F4", x"91", x"FE",
x"20", x"A0", x"E8", x"F0", x"F6", x"20", x"8B", x"E8",
x"20", x"C3", x"E8", x"B0", x"EF", x"60", x"38", x"60",
x"20", x"75", x"E8", x"B0", x"1C", x"A0", x"00", x"20",
x"46", x"E8", x"90", x"09", x"C9", x"27", x"D0", x"EE",
x"BD", x"80", x"02", x"AA", x"8A", x"91", x"FE", x"AA",
x"20", x"F3", x"E8", x"20", x"8B", x"E8", x"90", x"F4",
x"18", x"60", x"20", x"7D", x"E8", x"A0", x"00", x"F0",
x"0D", x"BD", x"80", x"02", x"91", x"FE", x"D1", x"FE",
x"38", x"D0", x"2F", x"20", x"8B", x"E8", x"20", x"F6",
x"E7", x"20", x"17", x"E8", x"B1", x"FE", x"20", x"00",
x"E8", x"20", x"DC", x"E7", x"20", x"57", x"E6", x"A2",
x"00", x"20", x"46", x"E8", x"90", x"DE", x"C9", x"0D",
x"F0", x"E1", x"C9", x"27", x"F0", x"D3", x"C9", x"2D",
x"18", x"D0", x"07", x"20", x"E5", x"E8", x"18", x"90",
x"D5", x"18", x"60", x"20", x"7D", x"E8", x"20", x"F6",
x"E7", x"20", x"17", x"E8", x"20", x"57", x"E6", x"A2",
x"00", x"20", x"33", x"E6", x"20", x"C2", x"EB", x"90",
x"ED", x"60", x"A9", x"FD", x"85", x"FC", x"A0", x"04",
x"BD", x"80", x"02", x"E8", x"0A", x"0A", x"0A", x"0A",
x"66", x"F5", x"66", x"F4", x"88", x"10", x"F8", x"E6",
x"FC", x"30", x"EB", x"F0", x"F2", x"20", x"33", x"E6",
x"A9", x"80", x"D0", x"02", x"05", x"F8", x"85", x"F8",
x"20", x"40", x"E8", x"90", x"18", x"C9", x"23", x"D0",
x"04", x"A9", x"40", x"D0", x"EF", x"C9", x"28", x"D0",
x"04", x"A9", x"10", x"D0", x"E7", x"C9", x"27", x"D0",
x"30", x"BD", x"80", x"02", x"E8", x"85", x"E4", x"E6",
x"F8", x"20", x"40", x"E8", x"B0", x"07", x"85", x"E5",
x"E6", x"F8", x"20", x"40", x"E8", x"C9", x"21", x"D0",
x"08", x"A9", x"08", x"05", x"F8", x"85", x"F8", x"D0",
x"10", x"C9", x"22", x"D0", x"04", x"A9", x"04", x"D0",
x"F2", x"C9", x"2C", x"F0", x"E5", x"C9", x"29", x"F0",
x"E1", x"A2", x"D0", x"CA", x"F0", x"43", x"BD", x"00",
x"EA", x"30", x"F8", x"C5", x"F5", x"D0", x"F4", x"BD",
x"30", x"E9", x"C5", x"F4", x"D0", x"ED", x"E8", x"BD",
x"00", x"EA", x"10", x"2D", x"C5", x"F8", x"F0", x"10",
x"29", x"20", x"F0", x"F2", x"A5", x"E5", x"38", x"E9",
x"02", x"38", x"E5", x"FE", x"85", x"E4", x"A9", x"01",
x"29", x"03", x"48", x"A0", x"00", x"BD", x"30", x"E9",
x"91", x"FE", x"68", x"AA", x"18", x"20", x"8B", x"E8",
x"CA", x"30", x"07", x"B5", x"E4", x"91", x"FE", x"90",
x"F4", x"38", x"60", x"FF", x"FF", x"FF", x"FF", x"FF",
x"20", x"75", x"E8", x"90", x"14", x"A2", x"1C", x"8A",
x"48", x"20", x"F6", x"E7", x"20", x"A9", x"EC", x"20",
x"8B", x"E8", x"68", x"AA", x"CA", x"D0", x"F0", x"18",
x"60", x"20", x"F6", x"E7", x"20", x"A9", x"EC", x"20",
x"F3", x"E8", x"20", x"8B", x"E8", x"90", x"F2", x"18",
x"60", x"20", x"17", x"E8", x"A0", x"00", x"B1", x"FE",
x"A0", x"80", x"84", x"F8", x"A2", x"D0", x"CA", x"F0",
x"0D", x"DD", x"30", x"E9", x"D0", x"F8", x"BC", x"00",
x"EA", x"10", x"F3", x"84", x"F8", x"CA", x"BD", x"00",
x"EA", x"30", x"FA", x"85", x"F5", x"BD", x"30", x"E9",
x"85", x"F4", x"98", x"29", x"03", x"AA", x"A0", x"FF",
x"C8", x"B1", x"FE", x"20", x"00", x"E8", x"CA", x"10",
x"F7", x"C8", x"20", x"E4", x"E7", x"C0", x"04", x"D0",
x"F8", x"88", x"A2", x"05", x"A9", x"02", x"46", x"F5",
x"66", x"F4", x"2A", x"CA", x"D0", x"F8", x"20", x"F1",
x"FF", x"88", x"D0", x"EE", x"20", x"DC", x"E7", x"A5",
x"F8", x"0A", x"F0", x"A3", x"10", x"04", x"A9", x"23",
x"D0", x"08", x"29", x"20", x"F0", x"02", x"A9", x"08",
x"09", x"20", x"20", x"F1", x"FF", x"A5", x"F8", x"C9",
x"A1", x"D0", x"1D", x"20", x"8B", x"E8", x"B1", x"FE",
x"A8", x"38", x"65", x"FE", x"48", x"A6", x"FF", x"98",
x"10", x"03", x"B0", x"04", x"CA", x"90", x"01", x"E8",
x"8A", x"20", x"03", x"E8", x"68", x"4C", x"03", x"E8",
x"29", x"03", x"A8", x"B1", x"FE", x"20", x"03", x"E8",
x"20", x"8B", x"E8", x"88", x"88", x"F0", x"F4", x"A2",
x"58", x"A5", x"F8", x"29", x"1C", x"F0", x"22", x"0A",
x"0A", x"0A", x"0A", x"F0", x"0B", x"B0", x"04", x"10",
x"0E", x"30", x"0D", x"10", x"07", x"20", x"68", x"ED",
x"A9", x"29", x"D0", x"0A", x"20", x"60", x"ED", x"E8",
x"A9", x"2C", x"20", x"F1", x"FF", x"8A", x"4C", x"F1",
x"FF", x"18", x"60", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"A5", x"7B", x"85", x"FE", x"A5", x"7C", x"85", x"FF",
x"A9", x"00", x"85", x"F4", x"A9", x"04", x"85", x"F5",
x"20", x"B5", x"E8", x"E6", x"FE", x"E6", x"FF", x"A9",
x"60", x"A2", x"00", x"A0", x"14", x"20", x"B7", x"E7",
x"8D", x"00", x"88", x"CA", x"D0", x"F5", x"A8", x"88",
x"98", x"D0", x"F0", x"A0", x"08", x"20", x"DC", x"ED",
x"A5", x"FE", x"20", x"D8", x"ED", x"A5", x"FF", x"20",
x"D8", x"ED", x"20", x"D7", x"ED", x"20", x"D7", x"ED",
x"B1", x"F4", x"A2", x"07", x"A0", x"07", x"20", x"DC",
x"ED", x"E6", x"F4", x"D0", x"02", x"E6", x"F5", x"C6",
x"FE", x"D0", x"EA", x"C6", x"FF", x"D0", x"E9", x"60",
x"A2", x"07", x"A0", x"09", x"20", x"B7", x"E7", x"6A",
x"B0", x"05", x"8D", x"00", x"88", x"90", x"0D", x"A0",
x"0A", x"20", x"B7", x"E7", x"8D", x"00", x"88", x"A0",
x"09", x"20", x"B7", x"E7", x"A0", x"0A", x"20", x"B7",
x"E7", x"8D", x"00", x"88", x"CA", x"10", x"DB", x"60",
x"E8", x"F0", x"05", x"2C", x"FF", x"87", x"70", x"F8",
x"60", x"E8", x"F0", x"05", x"2C", x"FF", x"87", x"50",
x"F8", x"60", x"A0", x"08", x"20", x"1C", x"EE", x"6A",
x"88", x"D0", x"F9", x"60", x"A2", x"00", x"2C", x"FF",
x"87", x"50", x"08", x"20", x"00", x"EE", x"20", x"09",
x"EE", x"70", x"06", x"20", x"09", x"EE", x"20", x"00",
x"EE", x"E0", x"33", x"60", x"A2", x"00", x"2C", x"FF",
x"87", x"50", x"06", x"20", x"00", x"EE", x"E0", x"19",
x"60", x"20", x"09", x"EE", x"E0", x"19", x"60", x"20",
x"34", x"EE", x"90", x"FB", x"E0", x"33", x"B0", x"F7",
x"A0", x"0A", x"20", x"34", x"EE", x"90", x"F0", x"88",
x"D0", x"F8", x"20", x"34", x"EE", x"B0", x"FB", x"20",
x"34", x"EE", x"B0", x"E3", x"60", x"A0", x"FF", x"A9",
x"03", x"84", x"7B", x"85", x"7C", x"20", x"47", x"EE",
x"20", x"12", x"EE", x"85", x"FE", x"20", x"12", x"EE",
x"85", x"FF", x"20", x"12", x"EE", x"E6", x"7B", x"D0",
x"02", x"E6", x"7C", x"91", x"7B", x"C6", x"FE", x"D0",
x"F1", x"C6", x"FF", x"D0", x"ED", x"60", x"C9", x"10",
x"90", x"07", x"29", x"0F", x"09", x"70", x"85", x"E1",
x"60", x"09", x"60", x"85", x"E1", x"60", x"C9", x"10",
x"B0", x"07", x"29", x"0F", x"09", x"60", x"85", x"E7",
x"60", x"29", x"0F", x"09", x"70", x"85", x"E7", x"60",
x"C9", x"05", x"F0", x"19", x"C9", x"14", x"F0", x"18",
x"C9", x"02", x"F0", x"17", x"C9", x"15", x"F0", x"1B",
x"C9", x"16", x"F0", x"1F", x"EA", x"EA", x"EA", x"EA",
x"EA", x"EA", x"4C", x"F8", x"E3", x"4C", x"AA", x"E3",
x"4C", x"00", x"F0", x"A9", x"FF", x"8D", x"10", x"02",
x"4C", x"D8", x"E3", x"A9", x"00", x"8D", x"10", x"02",
x"4C", x"D8", x"E3", x"20", x"3E", x"E7", x"4C", x"D8",
x"E3", x"48", x"8A", x"48", x"98", x"48", x"2C", x"00",
x"80", x"10", x"FB", x"4C", x"6F", x"E7", x"20", x"33",
x"E6", x"C9", x"34", x"B0", x"0F", x"C9", x"30", x"90",
x"0B", x"29", x"03", x"AA", x"BD", x"19", x"EF", x"8D",
x"13", x"02", x"18", x"60", x"A2", x"EE", x"BD", x"2D",
x"EE", x"20", x"62", x"E7", x"E8", x"D0", x"F7", x"18",
x"60", x"A8", x"54", x"2A", x"15", x"0A", x"4E", x"45",
x"50", x"52", x"41", x"56", x"49", x"4C", x"41", x"4E",
x"20", x"55", x"4E", x"4F", x"53", x"A9", x"60", x"85",
x"E1", x"A9", x"00", x"85", x"E0", x"A8", x"A9", x"00",
x"91", x"E0", x"E6", x"E0", x"D0", x"F8", x"E6", x"E1",
x"A5", x"E1", x"C9", x"80", x"D0", x"F0", x"A0", x"57",
x"A9", x"EF", x"20", x"3B", x"E6", x"A0", x"84", x"A9",
x"E6", x"20", x"3B", x"E6", x"4C", x"AA", x"FF", x"20",
x"20", x"20", x"20", x"20", x"20", x"2A", x"2A", x"2A",
x"20", x"4F", x"20", x"52", x"20", x"41", x"20", x"4F",
x"20", x"2A", x"2A", x"2A", x"04", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"A9", x"00", x"85", x"E0", x"85", x"E3", x"AA", x"A8",
x"A9", x"E0", x"85", x"E1", x"A5", x"E7", x"85", x"EF",
x"EA", x"A5", x"E9", x"85", x"EE", x"B1", x"EE", x"85",
x"E2", x"A5", x"EE", x"18", x"69", x"20", x"85", x"EE",
x"E8", x"20", x"49", x"F0", x"A5", x"E1", x"C9", x"E3",
x"B0", x"73", x"E0", x"07", x"90", x"E7", x"A5", x"E0",
x"29", x"F8", x"85", x"E0", x"A2", x"00", x"E6", x"E3",
x"A5", x"E3", x"C9", x"02", x"90", x"D3", x"EA", x"EA",
x"20", x"6A", x"F0", x"20", x"62", x"E7", x"4C", x"D8",
x"E3", x"A5", x"E2", x"D1", x"E0", x"F0", x"14", x"18",
x"A5", x"E0", x"69", x"08", x"85", x"E0", x"90", x"02",
x"E6", x"E1", x"A5", x"E1", x"C9", x"E3", x"B0", x"09",
x"4C", x"49", x"F0", x"E6", x"E0", x"D0", x"02", x"E6",
x"E1", x"60", x"A5", x"E1", x"29", x"0F", x"0A", x"0A",
x"0A", x"0A", x"0A", x"18", x"69", x"20", x"85", x"E2",
x"A5", x"E0", x"29", x"F8", x"6A", x"6A", x"6A", x"65",
x"E2", x"85", x"E2", x"60", x"D1", x"E0", x"F0", x"0E",
x"18", x"A5", x"E0", x"69", x"08", x"85", x"E0", x"90",
x"02", x"E6", x"E1", x"4C", x"82", x"F0", x"E6", x"E0",
x"D0", x"02", x"E6", x"E1", x"60", x"A9", x"20", x"85",
x"E2", x"4C", x"43", x"F0", x"0A", x"0D", x"53", x"4E",
x"49", x"4D", x"41", x"4E", x"4A", x"45", x"20", x"3F",
x"04", x"24", x"0A", x"0D", x"52", x"45", x"50", x"52",
x"4F", x"44", x"55", x"4B", x"43", x"49", x"4A", x"41",
x"20", x"3F", x"04", x"0A", x"0D", x"4E", x"45", x"50",
x"52", x"41", x"56", x"49", x"4C", x"41", x"4E", x"20",
x"55", x"4E", x"4F", x"53", x"0A", x"0D", x"04", x"24",
x"A5", x"7B", x"85", x"FE", x"A5", x"7C", x"85", x"FF",
x"A9", x"00", x"85", x"F4", x"A9", x"04", x"85", x"F5",
x"4C", x"58", x"F1", x"A9", x"F0", x"A0", x"C3", x"20",
x"3B", x"E6", x"4C", x"74", x"C2", x"A2", x"FF", x"E8",
x"B5", x"13", x"9D", x"80", x"02", x"D0", x"F8", x"A2",
x"01", x"20", x"33", x"E6", x"E0", x"1A", x"B0", x"E3",
x"C9", x"22", x"D0", x"DF", x"A0", x"00", x"BD", x"81",
x"02", x"E8", x"99", x"00", x"03", x"C8", x"C0", x"0F",
x"B0", x"D1", x"C9", x"22", x"D0", x"F0", x"A9", x"00",
x"99", x"FF", x"02", x"E8", x"20", x"33", x"E6", x"BD",
x"80", x"02", x"F0", x"AC", x"20", x"5B", x"E8", x"B0",
x"BA", x"A5", x"F7", x"85", x"F5", x"A5", x"F6", x"85",
x"F4", x"20", x"33", x"E6", x"C9", x"2C", x"D0", x"AB",
x"20", x"33", x"E6", x"E8", x"20", x"5B", x"E8", x"B0",
x"A2", x"A5", x"F7", x"85", x"FF", x"A5", x"F6", x"85",
x"FE", x"20", x"33", x"E6", x"C9", x"00", x"D0", x"93",
x"A0", x"10", x"A9", x"FF", x"99", x"80", x"02", x"88",
x"D0", x"F8", x"A9", x"F0", x"A0", x"A4", x"20", x"3B",
x"E6", x"20", x"00", x"E5", x"A5", x"FC", x"C9", x"0D",
x"D0", x"F7", x"A9", x"10", x"A2", x"00", x"A0", x"14",
x"20", x"B7", x"E7", x"8D", x"00", x"88", x"CA", x"D0",
x"F5", x"A8", x"88", x"98", x"D0", x"F0", x"A0", x"08",
x"20", x"DC", x"ED", x"A0", x"10", x"20", x"D7", x"ED",
x"88", x"98", x"48", x"B9", x"00", x"EA", x"A2", x"07",
x"A0", x"07", x"20", x"DC", x"ED", x"EA", x"68", x"A8",
x"D0", x"EB", x"20", x"D7", x"ED", x"A0", x"FF", x"20",
x"D7", x"ED", x"C8", x"98", x"48", x"B9", x"00", x"03",
x"A2", x"07", x"A0", x"07", x"20", x"DC", x"ED", x"68",
x"A8", x"B9", x"00", x"03", x"D0", x"E9", x"20", x"D7",
x"ED", x"A5", x"F4", x"20", x"D8", x"ED", x"A5", x"F5",
x"20", x"D8", x"ED", x"A5", x"FE", x"20", x"D8", x"ED",
x"A5", x"FF", x"20", x"D8", x"ED", x"20", x"B5", x"E8",
x"A5", x"FE", x"20", x"D8", x"ED", x"A5", x"FF", x"20",
x"D8", x"ED", x"E6", x"FE", x"E6", x"FF", x"A9", x"05",
x"20", x"99", x"ED", x"4C", x"74", x"C2", x"4C", x"74",
x"C2", x"20", x"B0", x"E5", x"90", x"02", x"F0", x"F6",
x"A0", x"20", x"20", x"1C", x"EE", x"90", x"F2", x"88",
x"D0", x"F8", x"60", x"4C", x"DE", x"F2", x"A9", x"F0",
x"A0", x"C3", x"20", x"3B", x"E6", x"4C", x"74", x"C2",
x"A9", x"F0", x"A0", x"B2", x"20", x"3B", x"E6", x"20",
x"00", x"E5", x"A5", x"FC", x"C9", x"0D", x"D0", x"F7",
x"20", x"F6", x"E7", x"20", x"F6", x"E7", x"60", x"A5",
x"14", x"C9", x"43", x"D0", x"D6", x"A2", x"FF", x"E8",
x"B5", x"13", x"9D", x"80", x"02", x"D0", x"F8", x"A2",
x"02", x"20", x"33", x"E6", x"BD", x"80", x"02", x"D0",
x"C5", x"20", x"10", x"F2", x"20", x"F1", x"F1", x"20",
x"47", x"EE", x"A0", x"10", x"88", x"98", x"48", x"20",
x"12", x"EE", x"85", x"F4", x"68", x"A8", x"B9", x"00",
x"EA", x"EA", x"EA", x"EA", x"C5", x"F4", x"D0", x"E4",
x"88", x"D0", x"EA", x"A9", x"20", x"A0", x"03", x"85",
x"E0", x"84", x"E1", x"20", x"12", x"EE", x"20", x"12",
x"EE", x"91", x"E0", x"C9", x"00", x"F0", x"04", x"E6",
x"E0", x"D0", x"F3", x"20", x"12", x"EE", x"85", x"F4",
x"20", x"12", x"EE", x"85", x"F5", x"20", x"12", x"EE",
x"85", x"FE", x"20", x"12", x"EE", x"85", x"FF", x"20",
x"12", x"EE", x"85", x"E0", x"20", x"12", x"EE", x"85",
x"E1", x"A0", x"FF", x"C8", x"B9", x"20", x"03", x"20",
x"F1", x"FF", x"C9", x"00", x"D0", x"F5", x"A9", x"20",
x"20", x"F1", x"FF", x"C8", x"C0", x"0F", x"D0", x"F6",
x"A5", x"F5", x"20", x"03", x"E8", x"A5", x"F4", x"20",
x"03", x"E8", x"A5", x"FF", x"20", x"00", x"E8", x"A5",
x"FE", x"20", x"03", x"E8", x"A5", x"E1", x"20", x"00",
x"E8", x"A5", x"E0", x"20", x"03", x"E8", x"20", x"F6",
x"E7", x"4C", x"44", x"F2", x"A9", x"FF", x"85", x"F8",
x"4C", x"75", x"F3", x"4C", x"06", x"F2", x"A2", x"FF",
x"E8", x"B5", x"13", x"9D", x"80", x"02", x"D0", x"F8",
x"A2", x"01", x"20", x"33", x"E6", x"E0", x"1A", x"B0",
x"EA", x"C9", x"22", x"D0", x"E6", x"A0", x"00", x"BD",
x"81", x"02", x"E8", x"99", x"00", x"03", x"C8", x"C0",
x"0F", x"B0", x"D8", x"C9", x"22", x"D0", x"F0", x"A9",
x"00", x"99", x"FF", x"02", x"E8", x"20", x"33", x"E6",
x"BD", x"80", x"02", x"F0", x"BF", x"20", x"5B", x"E8",
x"B0", x"C1", x"20", x"33", x"E6", x"C9", x"00", x"D0",
x"BA", x"20", x"10", x"F2", x"A9", x"00", x"85", x"F8",
x"A5", x"7B", x"48", x"A5", x"7C", x"48", x"20", x"78",
x"F3", x"A5", x"F7", x"85", x"F5", x"A5", x"F6", x"85",
x"F4", x"A5", x"F4", x"C9", x"00", x"F0", x"09", x"C6",
x"F4", x"A5", x"F4", x"85", x"7B", x"18", x"90", x"08",
x"C6", x"F4", x"A5", x"F4", x"85", x"7B", x"C6", x"F5",
x"A5", x"F5", x"85", x"7C", x"E6", x"E0", x"E6", x"E1",
x"A5", x"E0", x"85", x"FE", x"A5", x"E1", x"85", x"FF",
x"20", x"47", x"EE", x"20", x"12", x"EE", x"20", x"12",
x"EE", x"20", x"7A", x"EE", x"68", x"85", x"7C", x"68",
x"85", x"7B", x"4C", x"74", x"C2", x"20", x"10", x"F2",
x"20", x"F1", x"F1", x"20", x"47", x"EE", x"A0", x"10",
x"88", x"98", x"48", x"20", x"12", x"EE", x"85", x"F4",
x"68", x"A8", x"B9", x"00", x"EA", x"C5", x"F4", x"D0",
x"EA", x"88", x"D0", x"ED", x"A9", x"20", x"A0", x"03",
x"85", x"E0", x"84", x"E1", x"20", x"12", x"EE", x"20",
x"12", x"EE", x"91", x"E0", x"C9", x"00", x"F0", x"04",
x"E6", x"E0", x"D0", x"F3", x"20", x"12", x"EE", x"85",
x"F4", x"20", x"12", x"EE", x"85", x"F5", x"20", x"12",
x"EE", x"85", x"FE", x"20", x"12", x"EE", x"85", x"FF",
x"20", x"12", x"EE", x"85", x"E0", x"20", x"12", x"EE",
x"85", x"E1", x"A0", x"FF", x"C8", x"B9", x"00", x"03",
x"C9", x"00", x"F0", x"18", x"D9", x"20", x"03", x"F0",
x"F3", x"A0", x"FF", x"C8", x"B9", x"20", x"03", x"20",
x"F1", x"FF", x"C9", x"00", x"D0", x"F5", x"20", x"F6",
x"E7", x"4C", x"78", x"F3", x"A5", x"F8", x"30", x"0B",
x"A0", x"20", x"A9", x"FF", x"99", x"80", x"02", x"88",
x"D0", x"F8", x"60", x"A0", x"FF", x"A9", x"03", x"84",
x"7B", x"85", x"7C", x"E6", x"E0", x"E6", x"E1", x"A5",
x"E0", x"85", x"FE", x"A5", x"E1", x"85", x"FF", x"20",
x"47", x"EE", x"20", x"12", x"EE", x"20", x"12", x"EE",
x"20", x"7A", x"EE", x"A0", x"20", x"A9", x"FF", x"99",
x"80", x"02", x"88", x"D0", x"F8", x"A5", x"7B", x"85",
x"7D", x"85", x"7F", x"A5", x"7C", x"85", x"7E", x"85",
x"80", x"4C", x"74", x"C2", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FA", x"FF", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FC", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"A5", x"E3", x"49", x"FF", x"AA",
x"4A", x"4A", x"4A", x"20", x"8E", x"EE", x"EA", x"8A",
x"0A", x"0A", x"0A", x"0A", x"0A", x"85", x"E0", x"60",
x"FF", x"FF", x"FF", x"A5", x"E2", x"4A", x"4A", x"4A",
x"A8", x"60", x"01", x"02", x"04", x"08", x"10", x"20",
x"40", x"80", x"20", x"33", x"FE", x"20", x"4B", x"FE",
x"A5", x"E2", x"29", x"07", x"AA", x"BD", x"52", x"FE",
x"60", x"8A", x"48", x"98", x"48", x"20", x"5A", x"FE",
x"18", x"AE", x"0A", x"02", x"30", x"06", x"D0", x"08",
x"11", x"E0", x"90", x"08", x"51", x"E0", x"90", x"04",
x"49", x"FF", x"31", x"E0", x"91", x"E0", x"68", x"A8",
x"68", x"AA", x"60", x"8A", x"48", x"98", x"48", x"A2",
x"01", x"A5", x"E4", x"38", x"E5", x"E2", x"B0", x"06",
x"A2", x"FF", x"49", x"FF", x"69", x"01", x"85", x"F4",
x"85", x"F8", x"4A", x"69", x"00", x"85", x"F7", x"A0",
x"01", x"A5", x"E5", x"38", x"E5", x"E3", x"B0", x"06",
x"A0", x"FF", x"49", x"FF", x"69", x"01", x"85", x"F6",
x"C5", x"F4", x"B0", x"02", x"85", x"F8", x"4A", x"69",
x"00", x"85", x"F5", x"18", x"90", x"2C", x"A5", x"F5",
x"38", x"E5", x"F8", x"85", x"F5", x"90", x"03", x"D0",
x"0B", x"18", x"65", x"F6", x"85", x"F5", x"8A", x"18",
x"65", x"E2", x"85", x"E2", x"A5", x"F7", x"38", x"E5",
x"F8", x"85", x"F7", x"90", x"03", x"D0", x"0B", x"18",
x"65", x"F4", x"85", x"F7", x"98", x"18", x"65", x"E3",
x"85", x"E3", x"20", x"69", x"FE", x"A5", x"E2", x"C5",
x"E4", x"D0", x"CB", x"A5", x"E3", x"C5", x"E5", x"D0",
x"C5", x"68", x"A8", x"68", x"AA", x"60", x"8A", x"48",
x"98", x"48", x"A5", x"E2", x"85", x"E4", x"A5", x"E3",
x"85", x"E5", x"A9", x"00", x"85", x"F6", x"85", x"F7",
x"A9", x"FF", x"85", x"F4", x"A5", x"F8", x"85", x"F5",
x"A2", x"04", x"A0", x"24", x"A5", x"F7", x"0A", x"90",
x"03", x"E6", x"F5", x"18", x"E5", x"F4", x"49", x"FF",
x"85", x"F4", x"90", x"02", x"C6", x"F5", x"A5", x"F5",
x"0A", x"90", x"03", x"C6", x"F7", x"18", x"65", x"F6",
x"85", x"F6", x"90", x"02", x"E6", x"F7", x"A5", x"F5",
x"18", x"65", x"E4", x"85", x"E2", x"EA", x"EA", x"EA",
x"EA", x"A5", x"F7", x"18", x"65", x"E5", x"EA", x"EA",
x"EA", x"EA", x"85", x"E3", x"20", x"69", x"FE", x"88",
x"D0", x"C2", x"CA", x"D0", x"BF", x"A5", x"E4", x"85",
x"E2", x"A5", x"E5", x"85", x"E3", x"68", x"A8", x"68",
x"AA", x"60", x"48", x"8A", x"48", x"98", x"48", x"D8",
x"BA", x"BD", x"04", x"01", x"29", x"10", x"D0", x"06",
x"6C", x"1E", x"02", x"6C", x"20", x"02", x"6C", x"22",
x"02", x"78", x"D8", x"A2", x"F9", x"9A", x"A2", x"0F",
x"BD", x"8C", x"E6", x"95", x"E0", x"CA", x"10", x"F8",
x"A2", x"23", x"BD", x"9C", x"E6", x"9D", x"00", x"02",
x"CA", x"10", x"F7", x"4C", x"2D", x"EF", x"EA", x"4C",
x"4D", x"EF", x"20", x"57", x"E6", x"A2", x"00", x"20",
x"33", x"E6", x"E8", x"C9", x"0D", x"F0", x"F0", x"A0",
x"FF", x"C8", x"B9", x"00", x"E7", x"C9", x"FF", x"F0",
x"17", x"DD", x"7F", x"02", x"D0", x"F3", x"98", x"0A",
x"A8", x"B9", x"C8", x"E6", x"85", x"F6", x"B9", x"C9",
x"E6", x"85", x"F7", x"20", x"0B", x"E9", x"90", x"CF",
x"20", x"F4", x"E4", x"20", x"F6", x"E7", x"A9", x"3F",
x"20", x"F1", x"FF", x"38", x"B0", x"C1", x"FF", x"FF",
x"6C", x"FE", x"00", x"6C", x"14", x"02", x"6C", x"16",
x"02", x"6C", x"18", x"02", x"6C", x"1A", x"02", x"6C",
x"1C", x"02", x"83", x"FF", x"89", x"FF", x"72", x"FF"
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			data <= romData(conv_integer(addr));
		end if;
	end process;
end architecture;

